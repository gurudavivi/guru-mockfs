B�؄��L��X���s�pS[�X��<AHc�n��d���B>0*򕨞��=`���Q+d�����*���d�NՙC�ק!��W�^�u(�1��\������-���Vhݙ	�'̈́뎴�\��~�R��0���P��/Cp<��9�8��u�'2幱Ws xԘۿ���?��I9���s���M�]3����;삎���֡���	��� �*$ԗ��/=3�����S�/��-P�#���c䝲'�;��(�9�4�m�X�P����f��5	�o��?�0�5��6f�g��ʼ�3b^�K�{"�ز��
�J]M�R�Kha��:���Z�!�yPnˀ��Y'�.�)c�S89�r�x�������5,��JH���n8�5j�WW(�ݏ�昹�|XP�3�҄�ֺV����ί{i��Cd����Ƞ�ۃ��~�|�BS�
�x����Qg^5T�X��5�$�����sM��v�Cg��P���P�wn^xe�����C{�N �N�Ń�������<�C�z�B�O�T��O�X FF��!���dB����SE�G��ߎl���P]��5ٰ"��vS����q�K���@Z��N�����E�S�S#R��.�gI	�E����٥aYn�?���;��6`j�!����DdT�2��@6�������ut2��t��2v(��&�l¼Ң�B�N�#���8wо�0"���ǂ�hz@�^׳��I:�h��Ǡ7AH�k��a	R%  � �T�p���E=l���6�Z �ttE����S�����kX*����HXA�����06������2��~�ބӔiAXR�O�B�ǿ �l'	o����ܚs�ؓK�^cu�{���xV#�����L[<��+�:��Lh�����c�Y��'l��8]���@	��IǤԣ�����r[����9�'��𫖯�1�P"_lݴ\�8nK�2�a��0t*R��k�h&
D_cٱ��o����[ �"-��m(� A���L\���ܨM���G�f�q[ྨ���8w�x�V'P�R�D]�܇�q����&>a����6w���cQ�"ӡ��J� � ´�L(!E�� �r���7]�Ao��������V׎�� �%ɏ�B�9�^�I�mO�^�e��Ƃ�IO��qU![\�1P"0V#�zi0�h%��i��,S	<��P��>��k��"�q�	���\�~⫫�1x��3]Ko��Zv�?��D�g�)a�$�;�'�3������C�0L���6���Q�@�vT2q�{Q�pvE���n���0Й;J.�[]>fbY0��D�Bʹ�]����;��j%���_���{tz�YvAL�;l��pा?�Ʉ�B�c-,��I�yPyȅA�R������Xp�c��骓�G��2�W�JH}���ꈪ�i������2&RqV�ҎK��-W�.��-����g�,Kc�J��'Ʊx�]k�r�
�Zc!��
�ԖʍC��?��l���3�ҿ���iZ�`�,�ڱ��Osޔ �Ü6�e��i�pp q�_��\�AFf*�l(�-<TԌ�̫b�O�9rg��DF��]A�0/��AhH!�Q�'�k@�A�6\�SP\�hT(����� �ǫ^�k��}lcζ�.�b����RVV3J�B�)�o���eB���a��x�eҕX���c��U!$���O�bP��2����]�_���mA����#�=(D��0��������7X�k��50���u��3V�f:n(�5�q��.��=t(M�$��y���%ܨ�+�y|8��*���QI�|1�6��e���i>0hK|�_�(��S�1;�%���p��Yz-A<T�g��{�/���G��qo�t9�5bqcT��F�gv\��QI ��X4�
�E���{��B��� ?��-��|aل��+�?��r�
���Ӑ@�͏���6@VΩ�)�U����@�$z�!���������{+��ZJţ����k���q�y�PNv$2�����lFn*]�����B� �J�2U5���h�]�����~m���i,5L�l$�V�����7��EY5}�i4������>��7>l��ڕY&�
A����"�D��K�Zӛ*3[NoϪ�섧� ቉�0��J����1��Y�s=��mhq�%*gq�a��������4[����s*I�-���=���ۣ�}���ױ'[1�*���+����T�|@�:.��?�rΡ
W�%��wP����GK��1��k��B�����l�sp�Ao�<���(,ݲ�%V�:+�Bt ?񛋩�C�T3��s��)�nN�G��NE�?ׁl�V49�.�Aj������H6����s�LR3(�o��gՙ�wx��K�Q�^��*�8dY��bXHEB�	$�iQ�%�j�+N<���@�B[#�,�%]V�K�y 𦬫��<�g��8�'	����~A1��P����|� �<
%w���C�V[�x��h��m«,�A����l�mQ��C�240�O�@�s�N��}Ʀ�K�]�+ �d��:p���.�� -�5N��mE��.�zڇ�ґ�^[�5�[j�v�-���ԡ�M�1��� 5e��Kqy �6��bɈ}z��4	�N� ~��!W(ʬ�l܂P���mP6��8���S;�m3:�>�V�=ng ��ӞֲK�s"�P��ac��#�Y�^a�Б)�Ne���Qp�Sz�I�K��L������K�b���m*�V6�-�v} ���a�e��ϺW,j�6��'[-\2%��}�P��U(�i�Vﵫ#f��D��ܘF�&%VC�&����!��1�]��
j����5��D���(5���,R�v~���0���w8� �o���~:9�EL]ߘ[�/9�Y+�W�����-���+^SMX����,�T R����/;���'h9l;��]��)]V��T.�ϻ6I]e��Un}y�@���6�Y@w���-�Dʦ�F��O5�O0
���j�E�$K`��&�����kZ��d�B>�]��L:]��FT`Gmtj��s5�@J�Lp	-<,c��C�[�SE�`	��M� �	{���ٵC)(����G���G�k�������*��o�6Hw&k둵�Q�9�l�4�Я�X��`&g!��	DN>���[WIM�'�3Y3@��:��\��_�1i�$-��?7�J[� �);k�'�m�Lj!r�EثAY���u�Ȑ�a��~ab��g�5�P�nyl�B,�k���
��x�\��
a��;Y��ƽ5�J��JM� a�� ����c,�T�/�Q~��W��G�4r[��^��ˤ��B#J8�Qz�h#f!"�O�?I�L��	��OķF�of��-9
&N�U�MfxswE���wP�Њ�R�ĜF5��Dj��C�$x�r4�3��|b�1�}KW�/}j��ga���5��� ����"�~?,�F �J2֭�й+X8����d�L���2��d�O��(�I�܉�]���S!VM$�>��<<CjV�3G��V�k��n%S��]����}�̈́�(g�Rř2��b���Z�rBS�3�A�L��8|�6J���38�1U�QĮ!�B�)*Jq'K~w�vjO��F��(g��i��\h���
�q�]����x0b=��)��!w@Nv�@/`	�Wuv9M��S�RA�$��Pzap�:	�
���<[|�HtQ}��W��b�����ctKi�4����M݃J%NEޤv�g����;:���b�@���>������7�y��m�
�_ۛz�[�T�B��]�"|�j<���Tz�b<p�j���|n?w�ɀ:4�z�R�z�1t�
{�GN�ݶ2$~��[�)�UX�b�ww:Y0t�Zq#�Yt�j�i��> �z��-�S�H���U���}ό�A<!�~��%gcO�x�'��}jOZA<$�R�� ��e���l+}�i!I���s�(8�o[8�m&�W�T븀��cm�gCM(JP��BU�҅������Zs�Y�g�;�)6�<��LE=?���G�;�����]�Ͽ���UG���e�AR��8�J@o��g����K�x�uOk�O�T�
�tYYzG��T�]�~"/��FBƟ�t��2>�̫[Y_�+��⋓��.�p�ի5�ŗ�����ep��6ɍ���έ��f��2�f��
)�
��r0��r��1�;��=s�B?�j;s��H������cn.wlEC�>���} ��*�꪿{Lu���/��z�f�$D=���h��V�8=�O��y3ȁ`�h�����M.���O���P��ҧ�70�U����:2�s���"ьm/8tlAl�8=7��i��/���Ȃ���:
ԑz��S���u��I�q�ߝ�F�3����+�Ǉlz�F�j�Y�:��gVE��'&�w<����
�����U������*�Q+���\ˏq�:�D��0p_�I���O�������O�7�!�S�>
���o�s�Ǆ��+�G�dKJޱ��%ׇV�(��iW�v�OugV%J&����T*�hL_OR�;X;(u7]��1B���O���X4W]y�fB{�R'�(�/��$).�,L�C_��&%갥q.-�vE����꜕h#��3Gr���C��Ll�}�:�f�P��w����H񌱧%x[�H}Ts`v����kI+��(����|��p�i!�a����N��W~}���m�sE�.~�D��BE�q��8T�*�:�i�d��X�>I3M�}�巕�����'�����	R_�/k���Ж�{u'	��+{��9K�J���(�\
>���>ғ�����aَ<��ʪN;+���6eU� ���`���/	ւo���J��Uئ��.�Tߙ��ߨ�d��'LF/������J���|����,��Q� �v���	ӑ.����r��F<1�Eb�lG�V�
��8WC:�K�^j@���~H��ީ��`ZS�,�O���1v�9D+`�����AQ2L��1>��{��P�ƫcM˕��FXm+��ʏ��i��U�Yp��wc��_CJ�[TyI��$�i��$�)5�gN�41*-`�&��4U�f�d�E��o�b9!�R����ݸV5���'?��S�}��.S�����wՋ���_�y(D\�Mk�}��៶�Fwp:���=]B(0��&-<��hˢ�_�m��@*��D�}e����.f�����߾����P>R�54-S�g��V���YE$��;�W/[��h$ɐs{�?k�>j��|r?H��<	/D
����w���5�8����k<9�[HO�jy���h�}!u6��Y���HYEA&��*H�28����9k.v��0�t��6��>J࢚�0�Z��x���ד
�H�2��qܮR����uY�Z�*D��huɷ
����@,���p�A7hՎc@�6�m���ǁ�K�b�����E����ak@�]�o���S|r�P��&���QSV�3G�
ǭ}�KJ�yS�v!�4�����֭�&j�=_�\�n\�/���zV�SyL8N�S���5�<G���)d���Y~Eհ�SH4 �{�1Fc��ȇ
��*P�f�F�ۉ���0Ɣ�i��m 3>I7"��g!���HA��p=<�L�h"?:�w�F��ħ&�U`��Q�ܺ�΁�
�4�&�R�(b��^ߍ5�t؃�~�Ŧ?�}(#((�Z��8��O�j=<:OI��԰��հA�����DU����3V2vFSx�Jnó���ai���l�Br/�a�5��cI��`8VJ�á0ɡ�z�G�wн�[=�����b���bta�!>*v��^DX2Dv�͈ �� �K|���,ʦ���2GM't3tS��j��8��Vr���ݖ&�-"���seȕ�@�W�s �eư�9k�b�J�9Cik��?܈�Z�e\�D�a�"S|{K��&�~L,��]N�������2�_� Xv����s��*UD���N������v�$A�S��X��/H�6�Q�"�l���[�O�9�˗P�kI��h�8�âLNӁ��{�J�5]�}�"8�µe���lg6S�����Bu�Ӫ�8�^\j/u���z��5߲:��c8h�l�	�U���`)W���tr� ]i�\��V����LG��C�QB޽���;v9��#e¦8���85RP��S�A0��Pu��FP��J]�p���=���Ar����:Nufg�Y�/�F��ը+W� ���JK(��og\!��tXٰS;���
k��s�/��:\�{�����}��7F��8[6��?+�T�'��=���G7Ҙ��J��ߚ�<�'tΛ���ľ��k
`�w��y8�{k׃*r�D�w1�*����<i=o����GԼ�	Υt��<�l�#N�$���Bcr��_��i�΢�#���S-�%�ټ�-�ޫG�n>�Q���yG������e���>>Pv��u)A��z/��p��l��N��:�P��n���/�&��Z��F�SQyڠ�D�v�<�����]�.Z*�N]ȎP�J�$�����R�O��I��\�	����'v���M6/ $��|����H�뒵(�m!�%���<٢m��ʎ-8���h?j�r��Z_�+K�eحI��/>젣���p��9���X��N1�����k�l�R��E������Q nK���;�on�mF��� ��?���%XU�e�b��Br%+����ZfE�,� ث��(,Ʃ�n�"l�Y��T���}��(�:$׋�l���bc�j���Ea��WH���u����E��w���$Xs7�N(U}b��A�RL�R�(����TT,q�B�Q#�&�S�x�A��]���T��%�F�Ѭ��w��^u�:�B�����$Y��2��v:�JO���Q��<����!���L2�$^�����g8���hl�!�;>e.K�Wܜ�;Ί��3-�y[�5�63�H��]7�mg"�Ğ�R�%�g2ZL�	���6�"ue������%!�p�T��}�~Uen*v�h%q�ʖ:�t�v�|�>�g��ɠ�.A��� ��Y�@j8�ar�Ētx����_.��SPmV*.�7�:V�{=x�{��V%������-zt\X''#~�&
d ��=(t=!��M����?RB�%]��e��+��^)�OO��>V\^�E�}}�������y��P� ��~_������۔��fw|&��g��R)�g(�R�n��\0��]��)$c2'��XU8(j��oy+d|h��k��Β�m�.�4�B�T����q�,A������O�wWփ#�$�0P��n�\r
=0#��9�G~�I�[{�D��M�y����A�M��M����?��������	��Bf&<���N�q������8���(7P�D"Ջ:݄��D�f�q��)��rt�_ޡ��	2ew�x/�\p��>B���Y�D@����ۄg�Y0��[��s̯�	�=����*�h��߃p�a����4�ԗ͜\��F5��-��>I����_��;hP�_$9g\�>��d*gG��_��DG�Z����V�n���ͽ:p���QB 	q�aSG˙}H����	����?��w�;��V�ߒ�U����)�_<	�(dG����Y��׺^C��5�|�3��ϑ��9�n
�S����߀̗o1�b-�x^���8���5���M�z������
���XYp�nI��Y�r�א4d�p�S�q*������.+�Ci:������:F���"*c
��H$�m^��z�ܑ60�`,�h�J}��!�gJ��zأ�r��������:Q@�I�9���[�Z��eta��<��SD~m��[S�k��;�|>:5c�:�q������lA�p$���}	��4ݳ����W���Ngd�������?*�9���8���C!T�z�+z2�@���I��n���r��:�ن�Ո4�SV 8�@[
��[�?��Ƥ�X}� ����K����Ui�h�����r��uP��"%�]V�2��&�
u�'����+qR�q��	�f�ƣ��-���F�P��C��nn�2mI|�@���dǥ-	�T˧�}|����ݞ�b�9��s���ۦ����V?��SWi�DY㈙K:���M�����k6��(�rs���."ޜ`]��}���>mA-N�'�4�Kz� 4��j�y��D�"�RԆY2���FJ�+�������v0�-7?�?���5r� O�%Meta^\���%��IJ��1��rbn�H4�sW����)Y���E�|v~�����W��=C�d�%M���P@/��HTu&��W��*�Gp�� ��4�e��R؁µ�*�v'Y�^�!����cp2�@��)�*V�����4tj��� ��Y�~����쬷QHj�Kl�A"U��Y���2��V��P��m�)���M���jyd�ѥY]�=�m������	�S˲n��� �)���:�� g�]8���F�Ԕ_q��Q����M��o�����I�ŉ��wT�ϕQbޞ*�˥R{�n�dx\!\<8�:I���D�SP�����e�-W�\)��]#�"tp�� �0��s�"�� +�=�W�׽`�ڤ�ҶS4&�0 Z��uS �� .j��M���K]��m�啤lb%-�|򡖎�E��.xM��,���U-'
O�=�����̱�Ū�AL�n_��}��lnQ�q͸`�D�'�#�����v��
\�ۺ�0hg5��~y�0�|�c���¾8��ϓ!+���Wyf;}Fd�p
EWPf�>�P$�=���!:�yM���|[1�����v������S�A#� ��<Z)fɏ�3��2�Bl��?.���)�z�����15�خ�g.�A�l���D"�Ε�J7f�'}V���_`��~���WP`I�7��g�>-cܩL��a Y���P*3��fy�{���V��7Z R�}�(�_����5U�Z1�L�
>J6vv���gJ���/ɕ*3��$�>0��o+i҉�#$�l��QI}��e y���bSj�8��r�)�
��_�h���c~�4ܛ���4�<�@�1�5 �{��g���su2iՓ��t����+�#n�i��Q�3�(ȋ�����C�B�x�'����ܴ�0ɒ�m�[��|�ZY Q���b���	Jڣ���5�R R�݋�I`��ԧ4Mz�Ekkϛ�t�_��6���4<⹫����i(^��"���FԠi�q���5nJۨO���Z����__�v����ޤ&�i_�/�$gs��[G�,��=E@��6	�:/]`�-� V۳���v�
YYce�y���P&����]q���\�C�>�g?��uG%!���L"��uP�&\}̊�9GQpW�_5ccXp���|�0'���1�_�E{nbk�����џ�ƳN�	����"���q���0����~��� ����"�ƥI��X��T�^σ�(��I���ɠ3h;�юX�22��R�#>l�ԩ\[ ��J��J��fÒ�=��Co�'L����x�	8�3�b�!S��qN�@+$��(��Pg�����c�b(J��|lk���J?څ�� �0j��Q\��G
�$�
��' 2����[����r�0H"n*�I���Xָ��fFa���1�|���uF��F4��m�x�0��e��x�Vv�s���M��W�\��$Tf��!���?i�^q@օ���6FNX�E�֕���Fd��V���OxRv�q��Z�X�#O��	���r��	+Ke����?�l~m`Z��4��-��������?	Z+�%w��A4�L������]��پ��Tr������D���|�߯�j���+��k��E���q6�:W}��s!	�u�v�w�E�sI����K��
��F���^�3��eDU�gk�����R�����*0�ˎ�O���D�bD+����Oӄ�?D�qsdE�(��x��Ε���ܐA�os��(IS=e���a��~%[1_9�/�]���P��!D���e�6J�pd3�_���2=���_E[y/UA���1��T��\���t�:����G���5���*:�7c��	f���ֹ��	S��M�ro���V��o6�j~X�w��aD#a��3�gv��%xiY�4��n�~�L{U4�q��a����D
�.O^�=����0����֙��p��M|l.���*�?�r;���u���� 	��?X"��l }~��
��o?Aׁ���6�伫Bq�Xt�"������7���5����%F$�]�lm���8 Æ��ޖ�{g�H���ͺ�<M�U��	��}�m���	�M�+�Y�Ѣ�4�ОݜM"&�Epڟҙh_&�Tv��&E*��Hmו���L0����J��=��a�#Y�D_�^�uNp�N_�\%xCb�y� !�n\V�iFf���_�נ`�QP�*���Ny^�1'� [^K`�;U��)�� 9�����J��=V�(�r1:[����q�T�BrӦ]��PK�(Z�$���1v�X�$�g�h#��4+�!�{db�m���:C�+U�3����t'l��.�5?'qOGΧ?7�T"�lv����U����8kCՑ��u�o�E�@�y5S��c̓�g��[ʕ�GG+���U2�����綳T��]Z�b
s$����S��Ot%��X�|��s70-	�r^Z�\f�PS=�Ϡ����a�J�l�w2���F����Ds��>��4d���*]��*�8��Z{��eD��(xW���]o>y6S��~�����5�`k����M�]�=���J�e�Fq�v6��(�-�l�j`+QA��:��Ȭ�z�>���M�#���I�6��[�|��K�[��мNY�}]����e0 ����c{� ԅ*��9o`����Kz�7����#�86|���]3�v�l"�P�&��E`NdC��� �y$��l"��9����T�c��_����Eǭ���s�B$8����͂$���w ��W.QN�Ďd�_�X���XV���ޅ�B4v�t�#��9�FL�(f~�^�q"m�.zF�!d�W����� Dܨh�_��9���e�R1#z��Wa���`��'a�~�����vk�r]�dk�UƸ����M�c��ۅ��bl�_���2�����+qrC�1?|���&&�D�;���A	8�pb�P�\i�qlev�͛��✶���3/4=����e$�	�[ߚa��ȫ�x؛�^��4Pw��[�6�7�1�f���������4�k;�vx>h�]W�f0�oݕ�����I�8�����U�߶����!��o�N�F.�JGOF�m��ġ��@�7NK ��tW8,��⟀�M���x�&TjIY��D}��{ozd�3ڿo
8�Hǭ��r�V��w������L0���%�}��_������́e�{C3-����U��ٹ۸��ۅ��U�[�&ꢈo�~F�umW;���M�(���BUj����$K�w9`�?�J*��[�I?��SX�ʆn�2����3�J�4�x+�9|��~���ٷ�ǻY���y���Ҟ�RQ��N��3�t�Z�q�~eж��q�:r��m}��&R��*˲�=/ۯ$��G{3#4�JVV����%\�"��Jŗ�IE�[��MT�{+���y�A�.Ł��/��#�����CA��)��`���Hhõ��i={Q����#������D�&�p��E!�@�0��^(U��B�.^��0Ȍ��wj.�fҭ Bk>�	DK�(�5Uh�)�f��O�AIi_�5���B�TA��^cG2�y�VAx��XC�8�����6�S.��Ac	�pn#Bjm����sAǫ���p��>X�զ��z�re����bD�r�5~6[JV�-)Ⱥ�ɬ��Ȼ[�dN�n*k#�����s���M�-��(�}2�L��;�_�37���`x��|�TZ�#���6N1B�'���:R��`����Ebdf�@�:��]u}0݁ξcn�����.|��I�!�g�ܮ����etȎ�!K��9��Er�8A��)��6��q����ƣ��o��u�ْ)Z�!�{R������k��m��B�܄��T��ec�ͩ.$~���6�RY"��'�Jˌ�h�I��p�3}3�.jD;WV��C?W���_�e�e;J�R؂����(�Kz.��ki+Ku���]!BeV�
�;Ŝ�5�u��*�ܭ�e�@��xJ��u{��.�� "��.�٠�F�΀�w�9����w�R��u��1�XL2� �	��PI����\7��K$v��(}!�O�F��
6�%LT���d&�����D�������U�����ae�%�����Q��;���-O蛇ҳ�}�]�٥��%��-��0<PB����o���J<�xT����,�?�%�WS��Y翷v,�a%4@�8�~�G� �=�
g�T���˺�ץ��������{� j 7���hg��#�`��)�5���К��5F��=�bΆ�H�/�w/�_�.�u�NiZ�����,�7��V����qqDь`��Z0/.`X���]�,��I�i`�S�Bɀ��]�^�g0LЊ�j�V�Fh�z���(�����f.(�D{��W��H�w��E 𒇅�F�EɰnZg��}���d{v@���/�D�@Y$x"� +j�>"�9 N�C��x�l#���5���uZ��T���~)��SE(���	ӧ���j?(Z�'�c}��>J �露V}%�t;S����y��rQvͱ<*LR����(���O�0��{�ʙY�N��Ur\Ad�;U�Ġs�����3�)���z$�c�|߆�3�����"IKa��\�G������������'�nu|����!�oXlf��4C���k���C�b�fJ�V����C��؁����װ:ˠ*�f���
ύ��MG�n���ГB����S��wr�%"�K�[A>��?�2�G	y��0�D;��d<䧨���|�s5����.���M��i�U��L�8L-�H=6��~���7#�j�+'~�s��0�����R��'�I(<-syP�1-(�I�&pZ���vLm��HV��k�-����M�OOW�q�j�����i�����63����k-rN���`��������2� ��4����R�A����3�/$~6J4�p�l"��ܝ?��+�	U�2x��SC���%/��еX�<�ʓÈ���({@7�*֓bQ*k�/��$V}���`~p�|`������Cm;?�ٵ�����̥4��Ƹ��ു��}�N�V`g���v�\��^TO�<�E���)@y���5n�)Q��~�����Kz7�ѳ����9	��yF� ���݌�ML!��H#��G�>љ�bE�Вcb�&[\�K�,�t�ц(p�6��/'gG�ɮpe%Y�)���a�4��jlCA^�M��g�����3;�[������a����*��)�mDPPH���s'8�ત8Ә�	x�'!�ۢ]~m_���t���f��75��.|C/�ֽ.g���:���#���Ŝp�@�����J��e����<A�P�^�+��U���*}�o���Djʥ5��|u�4󦰴��e��!�=I��H��>��Bf;(���:�Z�n#g,*��P�%�wS/�\����JR�LW�<>�O�@�]�"IQ׭j2Y�<W�"��L��1�X�����4!�����_�4�U�E� ��3�d����V�P	�Zϩ���ljz"�՗�[�/�AQr������)TS��!�%�P���m�,>t�4	B�&����Yn��4���h��d�S؆��6ԛ�(b9���x��6Gga�������ܩ"}D���h�wfvD,����Z9u׸nJ�4�5!��52u@=�Qz��`��+,LD�*w�h�)�u�5DF��Ą�d��`�pX����I�^�-�M���WNZ���2��˕	X�%�ѾJ_���v��9Yn�K��-f���W~����m�7�3P�Q*�d��rW���A� ��m����؄,��,/���T	���PA�H��\�t�q/lc_+�/�.�/������M[�<̝��<����v�C%�e0A�A�������O	�H�6}��Cv褻v~s�>�	P�b�Tn��iׁwGy��ځ[�|J�>|Go͞��b{�Т��0 ��X/�ɑO4;a;$��J�v3�Aeb��i�U��.o��W9�IFP��`��5�os
���c��-+S;!�o�\��O@�?�
}�Ҿ�[�պ���Q3d�OղU���M��@]W{�qBf� Iכk<������C�V���@�Q�`�/C��#�:6�*E��K4^Ւ��y�I�L����Lʒum�#�d���[Hƀ��א�n�ObZ:Mkox�^D�k`N֨,,K �<��������3�.V��!�^k@k-^SO��PZ�P���uE��=5�����)=��TΑ�ODśTvϗ<�c�n/:���;�v���gjKK7�۬�O3l�1�L����Gp����f��p�U7cS�J�`�����~��_���������B�< ���� A�W^��P����yAf��?�o1?�$O!�r���IP>�l�QAF��/h_�ߍǭ rMz�D<�8�&=cZs�vv���MT�wN��([:s�=��X�,���>ӂ
)��3��a�Q���O����
p_4[_ǯ�A\��Ղ�8�*�����(T�O(�
�愭�n�5�b(��k���B[./{��[�$�Z�Hu}�Kw�+���_)�U�e-��u���K��g0��y���#�#��[�WПH�����r`ț�j��#1�� 1�0#x�����aU�h�6E��=�I�$@^���Jc��aTq��*���C�պ��\�_��/z��ɑ���B�R��YLl #dˣa����d:��U}�
�fԴ�>�DI��Y�R�b����ΊZ�?���Ihe�!�����5$P�7���+C1�yԤNkf�Ru�\18�4��=|�3wwE��^�\9�bR�N�����㠿h�y���}	���s�!Ld�Z/�� �L�~��|���z�S^b����Ky�/(��A�H���f�cS����[�OSQZLO��R{�n���i�W��SI��6��$:�#��sc����=�	b�䫲��t\8��}۴���`�pba�x˫�ss�<X@/�8�}��y��\�����)�f�cst��$�t��@v��#.��5y�����}��L�J��N�C����V���P4���י�;��AU��Dn�f�et/��ty���%+�@يQ(�њnH�v︧D�;���B���3>q� b��Ü�Ė�B��F��w_���33�_�"���G9A�?sگ�o���N_��-�?��KuY��K��d	�V����r�e�@	's�\�������T�)��xK����{]��¥r���iW�����Mu��$��5Ps�z�HY�k�N ��rՊF[c�T'|c�x�U��>,3�=1�m��{*����Z6�Z�H���V�:�6.
��(_ܼ8z��ߋЮ}6����B�D�+�z�U�p@"�ꇭ��?K�'�&�iu�󡼿k��s,��Ng�ښ\�VYxV'v���D�rgi��[n�΄���l���ɫQt�br۴�^b#Y
�]\^�G���R��w��+�M�MB�~����ȵ�=�+�T��-&_�5TT�<�]����UY�z*�پ>֢�����j`W�E�)��������-g�+ �O�!��2���!Q�3�Wxs�[Z���h�J�������`�M(�j�Zid��P�bf�|�la߮)c�̹rİo�媛�G���'�����xu��D'���픮$��v�G0k\�˚Wp�q���?��~B��~������GR�4s:�$�$������
�k�";��#��R,�R�W(�z�6u�H�I���ϥ�J��I�G+�so�ǜ6<����1�>���eI���&r���si��e�۽_ߧ�5�T:Q`7|_��Tt1�CF�|J�Q���vu���$m��eO~�K�&��aR�ƾ%&L�.s(�E��e�D�	��B)�ߵ�c��K#�ֆ�2�m^��}F�d����.���(�z���Sf.��t��w{o��+��r0���c0� ��3��B�f�e�jyw��;��x����������;����\�Xx�)Ҋ�l������ֻ���2U���x��b�p).�猶x���`���ڑ�k�O��Yf�����-�;��Ρ��Al����$AZ�+��f��ŵ��3�-gu�>T.�p�Ϳq�A��&��g))/���ݡ�>
V|�d�i=`�<
&��=���1�����Z������A�������=�s�̺�����PSQ;۷z�0N��m�3��m��v�d��B�aj��
�� O�e��fRڎ���"+�y�➘.B�����R>�Gh�:�l��9#��ܨPE�+c�,KɞP�wt���-Q�-��;���=���(��*I�#��#4q`���]���xo�h��e,ցO~�b@G�@{6���C�������"��H|a[�;����V0i�^��;#x��� \�!�.f'�I l ������h�7eڔS���.X+۞�i.�N��|�=,`ʖo�V?kz֪Ф;�����>@Q��W����<'��W��&,��q�bO�Խ^���ZM s���.���Λ?��ĝ�i\i)�qĎq��[��k��u*��扗��dqe*�d����/c�M�(5.��D��q��2�`�h:p����vE���I�s�$��WG���G0�������D�e���d�ɹ�Q�ɽ�o��映������ �޳R��nq��_iǗ�v���~�2�"���-l���H�WI����nB�S��T�^I�(�{B8x5q��e���z���	�2��#87 �
�y��HD�fw�}~���P�5
����{V�[�f��0�Z���-�|&{��u�c�]�?�f<}�����b���Dhڦ������Q�G�n;�RL������f����y8��T�jq�ƺQ�I��h��Z;����ٸ1l��e�D=Gqq�P��_""��3����A���� t�:�T�{�6�����%�|)�Z��$	��d)��	�F�=I[T ��p���{�X<լ;�k5Һ$h�#��\��OŻc������
���u�H�@e�g��m�U~�;鮜1�9� ��+>��
/�_��!��߫"����>F���#���h�ѡ��!�;�}$�9�ŀ�$���0[�Fhk��gM!4q����M����XPb�-����诬L��M�]Rư�J��&	W���:v�u�zT�N�,�{~���H�6�����&ɛz�^Li�"�ecAZ��R;]��q�#ꐞ/~O��d��hl0�� � 4�-�M�=CU/7ڭ?R�9 6���:u(*>���^����+F���_qm������f�u�v� 8�Ѩ��� �hN��E�T�����n�
��S?n�-��5���O'���{m�����?A�<ݮX)4�
W�	ԁ\�,%���]Zr��,s����>��cx)��L��W849�N%���]
q��Y g��,�xJ�g�38��q6�w�����q�[X��b,�t˩���|�!��I����}`|���8��
&S��},b��Dޚ5P����햱������gTM(��Ś$����̃�h�п!!�ʺ��-D֑�sD�q����v.�;����ʝ�,wck������~�� 3o�,��
�~~ٌ���9��JZֱ�Wd�~��%�X�@����nK}Ç����=Z&�q�>0s_zn��B�G����_���K�縦"h��Sa�~PB���o{�C�V�0Շ ��a���7�a9f9��o�C��t����I����Ps������Kƅ$�\�<$q�R�e��;��}�|�ZG�x������Y�pau�E浜�-������Z�t,(g�7�4��F���c�nC��yY�A���R�)���ߤ��!pҋC�4�m�
̶�T2���Vه��=�L�h�'���:��*�RE�#�@/��9c<w��<(࿓��0��wh!Y%�$�9��G��~z�D�(���?.�G,�\͆���0���%}0P���A�1B���EbTA�'$��Y�t�a�F�9�_C�ڰ��ۭQBA0U>�SGm��>�_w8����>E�����TN�Q���\o�;^�li%�_Y7m�(�A��|v�����K��p�T�~�҈]�jp�[�6��(zD`C[kWC��RNò��-OQD�۰�������[M]���.�l�@�@�RW������8Z��UE��==���砛E��x9�-�ދaX~�MG&��ȱ��i�^�&TZs=_�R'�cgm��vd7��Ge#}��-*ɘ�0�&���o��!�����i^��ω/;m 7�7,��G�c��!Z���`�2>��@��&����yN�޷�F���#�Q�%�t?_����!u;؄���%댂�<�r��$�w���ל0�\���<ی�[b"�A�ӫ:�"��,�� G��m,��=�����?Y���s����Q]b]bF	au��D[E�B����G�kͰ.t9zRH�^$n� �3�:�E�8��n���N���f4-[�o��Bsڡg��y����a���Ԥ0��Dn��=�t�I�>�f_�g0�+z�6d�op�U��T�8l������"F�������qe!�H��NI��_�q�ÎɁ�cd�R� �I0N�
�l�P�7�r���c�UQ���ݥ^-l����il��@L̐r%.b+�=<�j~g�����vh���'�Xp2:j�a�o���>��F܌-T��T�]H�1��˪��Ý$#?3�H�̒y��R^
n�[B��d�o%�>@9~C{^��%cnpNsX����9��v���ѡ`yP�c�s?��+8��� �g!ν<N  ޜz��,"/EkW��ϰ���t��6(	ba��O1����[Z8acn��d<�Y�;H��6>��V2�੭<{���d�'�.3�����CB�R�¨
�\���L��Z�䄑-�`�w���P����2��+մ6�*���$��KN���Kewb��v����t��H�����P,X��9X�����:�艸��'�2��[(��m�Q>�w|戆ٟF��ϒt�vo�R����Wꠒ�_t��t��v������o)aِ�����.B��z����Gu���
Х�_��>	�� ��Ԟ2e7qN�	�_���O�C�-�pFo�"��#��fl��Ϧ�ACb[F�!��\FI��ӂ�N*���!�`���a�ϋ)��?��3@���Ӣ F��Џ/]O��,�A*z/�,�C,�Q5h�$L�"[�NL�[���O��B9Fܻ�֙�96�FQ'

��	��w4��6�9C���j�(yS7�����$����Ɂ8ɫ�S	z� �����0F����-&+F �վ#�( !Lz<~��-��f $�x�U]���R�h��	B]��'�5�s��b�c|��������U��<�Cr0w�h@�du��d\=�,��'�J��vY�閰�6� �\�����@t�����z���P���*=dk�r�R�Gޝ$��r;����Y���:�>dp:��Ei�dFh�u�fįfOv���6)<�mE��#��y�(�
_QO8�Bぷ�3�{�3)���I6d!�|�V<�0����Lv2���lI�X|���+?9E�8�cz~����M��*�"Z�:GLt��L�%�(.���M!_��=�PQG�������<�<غ�3��2x�u���OYy���'�q%.����p�/e$ ��Y�ݨ�)�/ڷ%�;7�	�s]Q>�_v�Hq�B�M��T����MT�2lKQuk-��yx泋ܯĳq�u�o.r���~�Ăv��2�M�6-�\O�d*wZ2��X4ԅ7���c�@��4+����2/	fc��PP�4���S�@�P�e�7�5a�S=F�k��K�)I8J��-�?T؎���r�LU��;���Y�IU!+���Qf���f d��2���\-V���_�S%>�mC�;�����bs=���6L͐�0���Q����yFAU��F8��C�X�	=��/Q�YI�E������X�
?����
�qq�[��mB/"N'B�[yӪc	"J�F� �d�3�.�H���wu%����$��2 �>�4�����)2���rA7�@4c1�|;Tu�Ic�� �9�ܔ��b��y*�P����?��`z�5�QOT�r�}*-����[��(��w|y8J��'l�R�F.��pvE�s�;!��p�cY��;��ǲM�2�Jb�4m9�*hy2�A�	.�я6Ĭ������1��0��#�RR����e�Q���ɛv�q�r��"��e�o�_��t�5j6�e~M~藱_+�5���nxU�ؚ�=[�G���X�Vh,3_B2 Tv<��;�j3��e�g��)ר���sDw<dZzlN7U�s"��u�J�k�C�i���y�M��.��HΰF�޹c
k%P8�9d�-��])_'ee�1������4_�cd�2o_�g����^;0*yf2�-�e�@�r� ݩ{R�ZY)�%������L�)Q�K��Q�R��!���9Q?����pkˊ&��җfM�l��q���G�Դ�2����	����EO 	O��f���;g[0(�]n�r�?�Ü��d��Z�|`3#�R_�L���"��[fW 
ʬ�l-��-ۖV��y�#��uTg����6��5jĉ s	Y|�
���Qw�s��/G��y�>_տh�A��p�5���
�چ $�*�k�l�9m2٣ʫ�3ty/
2����H��k�#b/]awDnK*=�����P�`���~lP��'�:$8�����oyU?VX#�z������W�5�F8�Z ��
�*!�����C�cN(�B ��s���
���"�) 8Un�^��*JR��Ks�1~�ǧxJ��F�%�����Y��!u$D1o"�#ыKD��U\?f}6NBy$�}�q�&	�X�Ėp��A�t�U�VB��B]�k�:j�>�&��c�������(O�{D.P�Fx��/�z p�c�ߋ?ɥy@��y�X����N�wi�e��1�D�k��ˌ�,
���I�C�]�c��� � �΄�6�څ��Cy�����X�K�ضG��Dz��&j>�v�de-
�'�/�gJ���k��$Y�B�Op	E7@���#�hb�ULOk
 r1�ĂφN{3���?Y�w�$`~V8���0�8���R��-Kf�"%c}��刵@#�QBQ�զ�{y6��V��E�Ä�,���
��C`��Ѯ" �!2�h&ГuR���q�e� Ի�!84K�M-\uW�H��s����%��X7����>��sq��S�X�%F�	�XI*��[���G��_�)Ӏς�/� w�P�� �g��e��Jۯ@`�l�&R���&8؂$`�?����:˒OO;���Í)�-��mݯE��QC��.�[��lIi� �䃏�17�%�<�a��F|!����.S[�LX`t�շ7�xeK?M(���V���чe/5cRO�7�_�n��h^��j��B�|�+��
3E5�ZS܊Z^�"P�J6ӆ��"H�ZYl����DǪ/(��w��@D�2�D���>�~�������^��i%+�6.`u�H�h*��mc�?���"������J����x}�������VuL��CJ�b����R��+�g�#�����_�qb���HJ��0sK�*ϳ�;��j��;fL0#*Q���4)�d���ʂ�	�m��0�YH>`?�G��}����8�_SY�#������]uz�%�~�R���_9�-����e��Rṋ�z�\*4�P��7�t[�$pz�R�]�~]��x�抷��)"�*��c��P"��L��Z��s�m��G'�42�.&*EZ��E·���k=ã*;TҸ2�bE���Q=�G���{g�@��4��;\x|7]�mZ^��RT�M3��\@���Hή1��*D]�����0�yL���a"&]�Jj�UA@h��%�s'-^�m��!�5΍��Շ�9�?�V&�C{pê�%p����0�2�r�1bF���3G�Q�`.�hD���9��!sA�D�*3�'���r�"�;1�%RTj��9���h~�>��c*��N) ���e	�4�0m]`�#�H��EJ��<��6�|�LM�u�ٷ��γ��p'Fr��n�(k�a,�QgqO�yC4���b%=��p�|%'ub)6�j���1�{��z�`3��vK�D��.�*��	������
�hwB�2�-����i��܆�o+��99���%�����a�9�zבg�lR����ֶ�̐��Jal�L�FA%o1i��eq��*�ar�k-P��!���'�W&�H�
����Y�[�����#�٥�VFꟲaT^Π瘇D#�����X�d�gM�$�iV�S�9�5H�/�l�`WAlΙhw����MG������ʹ2�@9����qʓ�U��`������/�q>J���ϖ�G(��`����rO�����7�J�"��a���7�T�3Ԏ����`��Y���U@#��$������RY?�*��P&����/��u��d�/�d��Ēs_ocF3M	���k��]�a�_M�|��|��=���, +�wF�K�t�'�Ri����F:&{*ב�C���.J��#(-&en�Ҡh��s�����*xNB�!���e����<���ƶf�(H�(�.Ɏ.n�!�Xdn�w�+�G�J`5�EMZ����)�_�u���@D���22��9o��x�{/^�I��'˓V�T2y�gs�o��ЭG����7C_��$��T�L7��@~��ۗD�D!��t�z�@k�Cfd��\� �ۈ��}���2�I�).���o��F��}������W!�3����U��p��ۿ1�D��* v	�kSִ��܄�=�'�@"@Eej\<=#�;m���m�����F�fsm�[���/���MT2ύ�D��|�(�s�Z3qē=k[�Z��~S�G��PQ~�}�8c ]��3�>��+������i|�m[q�_��&��#*����kA�\���㢇����,,��<ޑ��*j�8�G#�����[u�o��;������Z�۶6蘹5���ySj�y��*���R��3*�K�_P北O���;�u��=z�Qw\ݲ���U=ψpGyN/�T���ϐi3� �}@˷։��U@M�qΩ8^�3�d�d��_�����Edި����~l~m�^����'㛅��F�۔����:wAc`s��>ۗ��`��`��%%�ZzNA�&��VR�w椡���u�B��"��BhޅZS?pQ$-^��7q��em�P��ʃ?�)��!"+bDb�0�j8�+���	��%�H�� ������G�W�)}_�j�kX�[�1J�Θt���ҍ�Ak�2+3���@��N泆{ĵ��%��Q_�(|J^���!3�=W��.U������\�:7W�x��9�*ܓ�\sS�wp�Tv�r $�8-bM�|���Gv�߉�x����b���� Y�mi601��f��R�����*XGy�{����R�O)@� ���F�?�]=����=\@��A?G�+�\콌~�O�E��j׈.m��b����·�����/�o�u�/j�M��X�lo����T"��1C�ҹ����M�����nq�Ԕ��=�b帷�z��@�,�����j��P�����{H��
�Ņ(��>������9��9H�1O��J����M��e� ����A>�G��#v�{�X��֌wGh'K@~��@���%2-xHd�8r�	���>`3�{8�	Vz]ur�m��[���#+�W[��B�o�@��f��PJ�Y��G��c#�iĦ,k�I0����Ÿ��%�3W�J�̮�� �^��9�|��c!���ϝT)��n�h9l꽬t�|�)��,+�愌Z�9�	}Gn�%嫢��&e��kaqhg4Y�A�$*���v�4�v&�7��ס�<k��Nق�bŠ�����$�# �����z����'-$��dgY�.��E*�����+��v�߆���@�ʎo'���R9#oUp��!�Of��qH�c��|$HG:��AF�v�c�5�Y��5�U7 �"���,/��gF�:��6��Sѝ����
��7hRYD�	�|�����kn��Z�1��x���~�d�j���{��(��R=��H%\���u���*k\��(�\��?�a�E�[�{�H=��0.������Ȩ�2һQ�H�.���X�SQ��� �#)Q��\&�O��O��H�6l+lJ�Fk��qb�rg�p�S�����RH
V�4x>��g.%'��蟨�F���?��~�0���G7%��eA�e�D�œ��$���>��wb~�۳)�u'�C��,���Ǌ��99�/s �zs�p�I�2o��2<~A4ؗG�(C���,�E�^�m�U� �*�ʲ��d��xL���(�C��Z��ȫI��߳���q�B~����=Y��&�:�Oe�� �-y �{�`_����}O����?Q�Zw}�Q-N��5�s��̼�4�mO/�d$��jS�Eew��4�C��5[.�:Λ�V3I�.�
�+l�AL�]��a`u��m��nL}oz��R�C�����ؓ�tS�5�t�Qx�dh-�m��8z:#2�:����� J�tP�А��Pԝo�DI��XU:%�V�_�����O�H+#���''���n>�=(OI��
��b��^�EzȾ�7����a�Q���ہ�������9G�߲_�pbm��$-vu���<oV�I��
���Sj2�h�O�̩B�ߢ8�[���Ry�H �^�N�?"�o�𼡉<MKˠ��rMܡ��)��ȸ�B�M��R^+����X/��\��^O:�6��Y��~�/C��נ�^�=�����^3�u[>�0ψG,bq�M";-����Q1:gr�W̪m��94�U���V�t�Ʒ��h����2�<X�uЫ�R��s�ra���!��#L�󞾳Hצ�#�#�b�]�����<Cm| /�E�X��=pf�����D^�'�o�w��=�cn�&��q8]F�T�s�B�wQ'F�pyr�?j-�RUv-J�,�v������[,��=�l~�1F'���t͹���4\3�c������g��>G).2v�H�z7��}��r6���Z�cP���C��l�o����`�v�^�9^5O����u{q��]�>��'�Q��a����sQe���C���냷6FB/��� ]l�.LG/�QIʆU�VS�� Bz�%e�{�ذɚ�(���9��OJZ���e.���0��:��m(��Uu 2# ���c�늗�Xʒ����Ij�|J��7�����fLPL\��~�2�ꁉ�➵� �Zj���Y�v70�dƈi����vU�7�@��H��Kӎk�aאƳ��{�n�
�/̷�-��l�o��I��et�^Є��+���߇^L7��#얦XA\�+�Vq�T��E�
��k�9�i�}.��.��gE/ӐGO�X�uRF� i��l�7�Q�;e�A;�u������ǋ�KX},��+�^Ż2�4ϡb�YmA�q���_�=6Ţ���iZ}8%�.��J�d`����nD�⍩�=" �������o�wό��:�f�
���w�<.��(���O|i <U�F�%���8����! ��d�P�Vkf��u�y�~S����p!��[pV�s�j��tA�\*��]H�/���z3M}p���gr�b,�aE���������Tۑq.���k�1;��
��y�oj�C��m��'z��O����=ĸH�r�2bo��~X,��$�!J�T��8l��1\�R�Ѭ�ϔL��uP:�(XϏ�Lgt���Bt���qv82�
]Ip�:D��,�\[P�]jw-~������9)���6�/p�N��;Dmؤ OA[,N�B�J���Ҹ%�u�x~����Ԧ������َ�^V ���5�l�U��Y�2������,�2L-���P�2�~E.9�� ��6�'O�h��H/��Ü�����2
�aοZΝ�� ��J�Ͻʿaڗ��RuU��AR�|R����Ls�[� 3������lu�������;0PU2�曋`:�L�6���eg=���k[��m�F~�EP��.�� /�{;��\�����92�TX�x���bN+����o�'�ʞ���rԍ>CW7E`H��V�D���RvLg��R�0�����⭝�V���(%q[�K(�f�>�v�"@T�W6�"��8V�d�ǥ����+}�'�4't\L�����O�7	'E(#��/+�n��	�OW�U�s���6�	F�"I�,P�_d��� uU�`�u1:J�<�O��?;.d3�:���'�J��a�����o���2��y��tfD��5T��hc�ן��=�$T�"JG�r|\��2��%y�Z�\�Y�z~�H>�TQ�J3]���^�!WPɡ���&�r�d;9��?m�DZ��/3�J�_E�ΐ��,7q#zdm���4m)"ú�=~��$�PQu���H۽��j]�|ȣܙ;9A��s6���]�*[�
�#z/���c�WEX{�w�e	��~�%�5��R�8�bgX�:��ְ)ȃ��ʖ�Oςs/�+ǯ�}���2#Ƕ��\�����{�)�/K�|�0t��n���3>@�T��PA�/C��B݄	���`�-�W�Ņ7�U�p0�X-�G��Ԑ��fq0l3�0��5P{��3E�չө﷐؋�漟�3�ܙQ�� U�|3!�P��)��CO^Wn3�9fM�wX�\��ՠu@��w���%)Z�zzp(_��9:1Q���Ux!˞L��a6x���D�Z��ϑ鵫�����O��S0<������y{z^�@s�b�ԤR�ĴL��rq.��|K��ϧ�<�:�A�˗�b<h�s�?�X��́Ji��� ��ۢ��!E=�%���kf:7��<qK�?�܈�Ƴ	tY�8�[y���qi�����q��:v�<wqJ�#��v����CEKu��\M��Q&l�#��4g����G�f�ƥ���g\�]s�%����YG��i�r>(8B�q��q$�h��A`�1��9�=}�"�z(yd�Q7�}q����X����NI��X��
,�b��Xo��؅��@���ڊ`6U�r����C��S�#�Ԯ�/���� O5������>�֦�V�L���:I��أ�Ox/ ����4��G�&�r͑�RS�H1�).{	7f(Z�/�n��+��S=aᆰ��1
X�����B�����(�J<p���9���\��PF;bC���2cR���Y�b�h.MٛM�%K�#����١��@��5(>�C1TV��F���D������ ����w����FPB�V�"7/hY�����0`����KWݑ�@��Q({À7����*O�S�@��\A�{�>{�^ϥN���@-�S�Q[���<��B@�`�R���$BU����Z���9�����*� �S'��rl���*8,a'DZ�)[!��^V_��`��=��X��	��8��6L��P-������(��n�w֕���t��o>[�Ko���P��=������B���F�>�*j���9����8�s�Mڷ6|'�ͺޭW�qB������J�^t��=Q��".����;�*Zc�b�C.��$����r�Y�M"8�Q� +�,���͂I��X�ր��%BC>�.{��X�2�+��9�4�9��-rF۶V��.�K(�b�+�l�#2h��i ���ޠ!��s@���p��ý��LƢ���q	*ɠ�a����Jҫ7��b�8��&e����kU~N��������]��@�"r ���6,go����+��/c/����'/g�kC&�:���c̗l3�a�6C�m���q(G�_����!`��� �ĄW�.�$W��b�9�܂�k��3J��׵^�r%X|h?��mI�o���Yh��/w�	ǮA0��\������PQ�,��Ҋ�Ÿ�/��Tc[�>Jg���s��J� x�$�N��,C����\ԧ����/u��+��[�O�d�2�r��y�(�x��~W���r$�눿A;�eYc��֛��J�]~g{cV�(�E��sϨКK�=���)nh� 0�D���»	���i�=�r�\��K.�;���0����<�>l�A�7��+���P�Q���t����е����F�,�B,�PHaK��p,8N7BD�"֨��4����=����ot%MQ��ه@�lC��gi��׀x��
��.e��Ĳ��܅Ų ��-X�Bg=��߹E8��z�Eꔭ��k#�
��;�3$��}c@�2�f��C��Q6�2�Ф��t���������>�]S���DQ7�V�k"`���>�(�qb~�LD�ֹ\[V�Q���2,�36㕩�vX"Yl�z�`[�׺�7*#߱���r�0[$U�+BP��B��V���h��2�I>��u�n����[�<2a����s�2h�4fY�T�r�g��"B�#0����A�O�Iz{��>���sc~QL�
��Y��g�'�GX8!��ez�GTVv�������O=�t¸�K�M��&��臬�jFi�]N���E���x[J�N7�!ߐ��U.����ETpwU��F�=S�c�S��W��:%i�"7��7!��,ۊƦ�`����i�+7UT���c�x4��`�H0g+��k�|pmP�aYp�N&�H��v��&
���M�"�(����*>�2�F���<�k��1k�qsn3�R���_0��"�1 d,�;c���1�uC�CFi�b;��Ch���}�$�@p�h�ۇ�k1 ���^w�%��4���I��E��=S�?Ο)��g�J ��սB���x�,(�~���͈�As�@v6u�H�O+�d@d�V��[T:�q
aֻ\>8/4���-���63�t�x���o5�ٳ��`����7�(����\�eZ�>�+u>o�������0*K\>\�"�<�qx�L�^�u�1�`48�;�#�֚�c�������.�c�� {@w���@T�����;}9D,kB8{�Nm������i�n�������M3#-T����FnΣ{7m�K����J�q����N�EA[
$�k;�D�[�޶e4�����QV��tk@���?$��9Q�B/��"e6^4Sfb�@����pa)�;��]�"������(�$���I ���Ψȧ'.�gc��7(ݲ���cݫl�OAzi���eU����^�����_�*��Й_h�E�h�C���h���z��:�ٷ5���/߲��yǀ��٢�e�k�Ԥ��D�=��G	t
��(��w���lϕ�8ƿ���ʊ�`� �F;�C�mb�^��e��%%��I��Z<d����8�o$8���|ɮ�v!G��ט�i�+�N�1g!@�`E�֍sO=P���=�����#CX.���]b���i�g�S�q����r엠�:�T��'2������Ϸ�H~��=��vx
�$��S��>��"%׺Y�@��.�t���]��JO�9�L���R[$ǘBH']!;'��ez��e�B	���0�:��hP��E�������{������5U�Y����2��ԺΠGhD�7#�YjV7W�n�1�e2q
���UY5�'�X�1�ch"ͨ�7+���S�����@04�A��Ӿ9Z���<q���>��#<�<��|m���W�B���_����1jps	(�Sa��5�<�6w�m��FĹ<��L�����	�G�_'�?*�ǳ���/ �A ���M����s��hn_��+N��[��_^��D�[�rܠ�L}�ft�+
��y���M��G�,
�\c~�Bk����P���[;����#�{ě��@$��=�JF%�����롛��M:�u<�cV�Y�/�\z`�ޕ.!�L,f5e��.�0��V
���Y�~Xzp:'���Ǐ����N�C��%��H��s�S�-��c�峇�kV ��ꮡ}�����!���6�4��{FT �N�A�ei����D_��\Z�?��I1\	gY�t�O��(���^nt6�(���=]Co�F�Qp��)[ԦL�`S��m��E��@����'�_W��0�k���*qzD�����%��(E�?�`�R�����,g�I�� ��I�'`(Џ��J� ��M�t�ֈ�ɕg�Ch�q˖|��2ͲOE1W�;��)������6��+NHZY26��b��ޅ]I��OQ�z!���T���aNJ�a�P�Y�6����BA<� �o�E��ECX�
�_0PX�❑�)p{�QC�ĺl��U���XU���60��q1���P�N#c����sM��WM ��^͌w:8c�
�ȉ�s��!߉Я��6��)4͖��<|$��@���u�W��
��j\��$O���z4yy��8�0 �F��&!�3z�zNr�� �ۤ�}T��l����Q��4X�{�̃N�Pf�4/�.|�y5�O�h����C����fOS'ϯ����G����r�/���ؾz^�ZD�%�! <BA�Y�a+!L��\k��(��< J�M+�����R��)��G�_˧��݈�)~A!w�m���nJ�
� 6[��D:`f˰x�(��|F�Nj���'� s��%3m�Mn;�y6�y� p��*�R�/�Q������J��U�S���#����ɕR7%
0��rjÝ�� Jh��1�V�V?W�����4���72j)�&�� o,|M�{���1��I�2��f']J���r�0tpL%�#��*�a�H��c���G���I�ndp�Ix`*̹�yU�x_�O���,JZ�OV�����l�������PP�x������Mx��)7τ̂��\ٳ?���.O��@�F��I�~|���M .���Ѿxց���PZ�y��6��s��:�Q:H����TJjE�m��Қ	�eah�ڡ�nn���1=cL�su{y�s
ϸ���F>e���.1�1�-�,~�Q�J�C� ���(;��\f[�ץ�ӀM;O�����Kw����δ|��Q���Sj>]O���J�܅Q+�3`I
:��֥�<GPSA�k�3C_��Տy!��]�^�1�쉲w�4l�e��	<�&�q�:�̔Hޭ��o����(�a&G2�k��y��b�s�S4}���.�,"%B�E���~��N�E��{zt5�K��"��Og���ۋ�G�غ)�Az(}�;#Ĝ�Iy�J���9��$X���'YG1�.Y{�O�ˠf2��y4/�h�2����^�rZ�v/Q[����a/�Az�9�2��t�-A<�#t�#���g^Ud�1���Zz��k �ɯ8�H�l���y`N^H{_L�ҡ@ʔ�p1ɩ���m�EH�Z������-!ۭp`���㖙/A4e��Ph�9��pre�]]	Wv���,!��N��h�&%qoĠ�����.�L	�T� �P���?�qrֿ�8��c�uv�Ձ)��L�1"y��4y$��n{� ���٢	��y盏���0�7G\|����!)8MJ[d��߉ 	lD�E�M���aj��i���0h����,b՗����8�v�M�;&Z�`@������8���ܴF�:�	P�3"²2���HƱE�/��W���]�aeL�=G3Z-��R��_�Z�=����������������A#�+���D��ўד