d�����~���:�#��,��ٕ���#�]D�P��]�od8{/�.	V�t�uL��F8\�܆���lܛ����R>ײ�"QG�R���e��>-����+�Ą�Z�� ��g|қ~�O6R����ݕ6KV���`�����1ۉA:�P#����nt�4T��;�p	����v�\s
B@��].iul:J[b��T��f�+P"'`�7�'gf����w	u���.���T�e���D,;"�h��E�BP�RƺL����nm��o�>�X��|d΁@��w��W�}V�"�݁YB��u�;� $V������ r[>5��i�H)�'�����e��פ�a�l����5���:��_'�t��۸�I�J疼!8�s���h~���w؏�؋᧌�s:f4�U���67��A�a��	��SΜ����B�U_�i-Юj���z��-{�T&)�dԕ
"���i��Zfi��Xw*�%��oe�-�G�FI�j�M���������j`aX�D�9y��v���.8F���]�|�y>��& 6i���`��&����[�^Ugv62dx@�/���rl�vׯ���G5�e�)!�֠��@��1�e�G^�h�>V�f'����P����I��[ǑQK���7��_/�����������P+��7�ojf]���`s�dk�d�o�cE�B_�j�ljri��a�"�e*�%����z���!\:k.V��_Bo����B�c�Q�ś/���i�aݼ���z��@��;PH�R�,�D{�֐ªd�;Z啳a��/��8l��J� X�2F֋yR�o/Z��,����bk��3��@I|J>Ui���5|50���:S-LGM����Ffڬ�
�uOTK�/��&f7l��A~���f�aA~	`_:�j��B�-�W'�.��G��0��K��ԫ`q���!��k6*9�-҂�zz�)k�M,��%&	�Rҝ1˫�����g-]�؏k���AS�߷僓�%gx����l8$9�2E��c��I��:*��i�nF�n�/��̵1�.���[lY�8/����|���@�`|�AT)�"P�����ջ�}����n�4���AS�'gDn��l����]����>�m0��i�X��"_\'�R:�:q�&	Ѭ���� tq;r��+p!����ѻ	�W"xF��H�޿gC72��`
-#-~|or���l���k�Wj���U�Ba���Q����QM�r���s�3��Ap�q?�!��y��#Ss�D�6��Cu�n�<�&H{��$��[��]fXrv�i,��4=�_�����a��ͫ陸���	�->�`�R,D&��Ӥ[���Q@k�}e�	��y�!�X�����-m�V �ɓt����K6�hp3��;lQ?y4�M
~�m���T����Ͽ��<`���%�.X����k�][������K�X�2U3����_�>�:�y������C����R���R�����������k��7F����N�*�i�ݿ �z3
Uɋ�C�r���M��K�H���f+R�A�;4l�0w�D�n���s��
JL����1'����Q���T�{�	�Zɤ��@EWQ�6Ԃ���"���10�$t��j
�f���=�Jn}0�)��Z`��=��d��F�\<c�y1DPǬeT����W��lM��	jF<�â����f�i��~wVd���Dc�V|U$��b1G��[q������I	"`�'�`�񰐆�F��J[��+[UX�"�U+5kWc��+(�⑤˶C�dbb�o��v1�&ƅ� )L�hS�?a��P��ο�q�������&����`!h�6�
�R���q�u��r�PR�,Q����z?Ka�|z�j�����<2��0l7�7[\AiiY��>[��#O�_pq�[�p䈉
��zh����v
��ˈ��~�}_�D	���9(=���
]i@-f��~{�.LL���g�2Olʕ��S>_L�e�k���~Ó����,�A��gOBE�>#O�͹ܬ����,E�w�:wa}J�����c؉V ly��1y,}t����d8]R�O���Y�L�I6�`py �Fa��25Ҋ|��`�N�J�adMK�\����1�u~O���ȋw��U�B�R�nCC%����k2�E��;��!�f����1�6<i�5�!�1K�Bu8w<�B�k���ם
~���;�ʍ��J��=\�e��]�����Y仌j�-@g��W�.z幼z=�_RK{r�=�� n�~p!�JS��j�O�rh��oS�(�����Um=3)A�ot�����=��'�-K�O�@�"�P�Vͣ�]A��-Q�f�����.K����n)%���?9�Sj�a�-�I��*�T��>�ٯ�܆^,��k�j��}N+*ߧ�y"6<�J���9����Z$�1�0,grڈ��������*�SM���Z(ͨB�@ڪ���<���x���cQ�٫���PP�e�k!��V��Pڛ^yM��b��v������SsPɀ�[��7��_|��,�|�}*�j;���U��<���ơ��(0و���������pk�.0U�����?:�5�J�9�&�p^��4���g�Sl��c�J�sA��~��z�j�l{�:�0+38�o��-a�ǻd-�>d㛅�"��e�b�"��qC��f��x�Q+�g	�`�}6= 8{حՑ7�q_��E��+�/}�6�i�@'�nS�g�o���h���:���g�s�4����w�Y�!�.�+���d��do��HU�4NIu���b5um���	ڜ $��.2`B���%J�Y����|W���n��(B�%��V�zߢ}C���cDHHc�F�nK���tI�G߷ǩ���Ӡ|X�IP_���b������hFY8c�`]��ا�R	zG�d�_t��q�'ֲ��V�Al`/���ʩ�o�L��K'8��<&-ɻ��,�����/D��-xzU~"�|JxM8
m�E�_l5�Q�6R5�n�EY��?�X�>��S�ްM{���4:��ό�]"T��)Tɗ�T��z��!�*��o�#����F��%���9��f������c�ª��J��'��r�ۨ�ʕGeA�P�O���*��Jv+	_~�����T�a��7Z��n�(���j 1+3K�n'�A;�r�#����ydɃp�i��K�T���Ɂ�I����1��ny�(��@)���U��$n�K#^OI�#J��H�bf&$�3z���J���Lo� �C�+4_�k]A�Dܷ;A��3*�Y�fP��W���:�\�כ�~�Z���G-G���e54 "L�I������kH��l��E(��?BU>��Y�O���LX]0�	���V�'ѭ�J\Yy �6W�f��G\}?���cț\7���p+���A��;�?PM֫�t���Z_.�*�������\,ʶ.���v�	����s�F���^����ό��Q�	C�"֥�X�RFJ%.��y�2U��R
, *���>�
R�u����a���P��
�T5+�x��yc�̚on\���Ig�|},��Ī3��z��?W�*t���R Le��kS�l��r�t�<��Er�1Æ;�m���7ඝ�W��p�$ت�z��M%�1�@��:R��9��49����'�co/je�xۡ 4Č��}ɷ{��/� �9N��f��k��#�4��#��rc�ՀP�^!g���;"�0�H0�޵�D�e�G��e���������uF�N~���8�	Y`xl������z�	H;���66e�c���m�.a�n�:����?��,�>w�41:e~Uߨƺu �'��o�b��!�W����/�Fm��<[���"FÝ�Ɲ��� io�4nP|@�Oi�%3V�����I4P�������cX�1�F�m�R�r�C����y@��k�#ď�\$7��&�+nZH�).`�����^�;�Y2}���_��:d����{8�����6���Zb�VA�[�/&XufyߟGc!���-]N����n����eu��}���N�b�l:,������_䢹��PX-����)�Yˍ��;>&�ߧ�]����'/�|K��v�~���X��h��f�1�tޖ�Hw���om#�B��J��U��4	�*�2��q�� �mԽ7�7���'Wmj�����Ǆ̬���K�`\�L������8ͅ"lI���צG����DH���
��F�+���F
����.<@���JZzR*>	e���g�x��K뮑�fյ����Ⱥ�1�*ӦdH�q�-�:�Ē/��s���܄ ��?��.ɟ)X��m^% ��欉g����5B�=J�`�I=���6F������a<��Zǌ��q�#����5�9�|�u�ti��.K��k�`e�My�t�P�B�s������x X� $�s~�)��ҍ�_�r�%��	f��!e�ᖹ)C�f`;"Z��6�v$bb�f���D`o�P�GR�qώ!��v�Ϭn�	ł0-BO�T*�
��,� ����=���p�\!�*��~
�\���9�����5Bq�����ڧ���lݰǞ&t�PI;�f71�U8{Zx���S��hE](.�=M�k�|�k�XJ�$��Y�MB��8P�I����v\�����1V�����������w|����o���Pr[{��v&���<�"��H�_��=�)�5Q"���ͤ�o�`�������`��S��q-|� ,�&C~[�������[>!���߲�3%����'������٬��f_-~.+f��v�)|�L�|�Jc3Pdn:
��ڌSK0Z�����S@��ի/�ш��xۿ���k|:��q�
Ӝ�z�x*������(@�Z�<�ߑ��\k�S��7
���bpP����V��uű P��\���T_�wx��J�"?z� �j-�(#�۬���D�}7�$~ި�AN�n���غ����h���$]��,��w�,�����������6H3Ε��2��c�����X��G׵bh���U����p��ƭde�ئ�%�j�"�����Ȅ��T��8"��B���Et�v1��H��»������WLr��ګ�r���X�4��������������<a��ͯ]9@`�-��H���7��c\J�i�s}w�PƻKi�e��E�T�53��_�x��#�O��҂�����2q)���� �v���||���?��z_��M���Zʔ��@	���GR<�H��v��?���G�����@���3�vȵ{\��)s�0�|.���E�x���o���U@LNQT��uhL�KmnE��`Jy���s ���U#�n!?-@�1\�
�P���|[����p;���빢C#���{u�w��P��1�,�7[���e�E�n�-��G��Hꦭ�ouս�����ޠX���KN,�yT�8@϶����r�Y5���1���d���H�U�M��ALt�+�)�]��}����_�ÅM�;4�}�+�W;9^(�u�,�ze�n�ɛ�h�,/3�S^dr��ǁ����%��p�f����?���ּ�}��i*۾g�*1�h��iن��T����Vu2��_k�W�j��:6GB,سz�Y� ("�H�k�_�Y�N:S���oX�o��'E_�M��"Q"J�[�>�u(�q8���G�G��x�i~X�fLhΒ��΢]��
@�I���1�JI��_��ū�~� �V\�9t���E(H[�1UF-�0l�f���lY�y���R�q �ՃŖ�_h�<�7���]o`�a�.e,�
c�ȰkC=�M���y�0�F��f�w�J�|��㆜��E�p&ڼ���F�C��O���k�G�O��@����)�N��v�J��LSڞ���h�+':i�}�T�8�!Qs��:Em��Ő9+�q`ΧU|�>0�}j�D��ϴ}�A��S���G���x�+E[@���%���a���~�B��6���5��+��7�?��w���&u����I��V�*���#S<k�>�j��NwS~�F�+�/o�:>`��^r�ڹ{La�R�C�<��q_x�%pd�?���Y�D�h:t}n�=O�>"���8ڋ�O����lD���蝖H$�o����d�)�@��U��EXJ��,�f��X����ì6��l��J�QGN�!B�c_���� �Hm��v�6��Ȧ;�-�~���$�ʵf�\�V���K�Ќr&�އ�8���FME���<���$��e9��;�Vf�	Q�6�t%����#� $E<pi�H�멗��� ��]!�i�7��(��XN��w��+�uU����woT��$�uY�l8�6��C�V��y��������]�|�(�~�G�M���D��~�(�t6��+~�6	MϮ���TI�H���I���"�3,����o�jK�a�-�BQY�.��О��S�Z��8B�;�� ��"��z~�i<��E���qZmZ�	��I��k��~}�&�a��眖���������8\5���������j�_�H��ў��/�ݤ�"2�j�W ���A���؆���u�(���E��ɶ�Be0(�ex�л^1Od~�a���0D�J���0Y�"�AP�r�%0g��"2�	�2�ճr������p7_+���5�n��H�n��E}GaǞ�#�Seq�n˰1M�n8dB�Y�̇�(�KG�pU�]J��Y<[?��ϩ̯p[��X���j.�Ox˃���'���C�	���2Q� p �����ގ��p�\�=���Nr��� #�q>O���r.�g��� #��Ϧ҂Ew����� ��6B���1�A����r&�SLX�?���%l��G�%PD �҅DD�}��z�&�T�ʞv�*|N]ݺ��6���lS�0�� n�z�e��)�R=+�����Ki��{Z�W�����\���ݝ{Sw2P���_�=y�@��B����:�{�Yd�@4%�-��F:�q�6�2~�F�1��qD{Q9k�սOjɋ�ՈRÑ�eǬt��;�\x��t���c��A��ƚr�J}��+)�Bh�B�\1㳴�%��Q���FMt(u�kH����=�#<`~3����T�����s�8{�O嫧K���ʯ��"�ˆ�}a��N�=�����чJ"H���&g�!j�S���R�14�K��V\e�R.�ym��Ǻ�4jn�������D����yRJ�]�.��/�$�V6�� Ϳ�b?&�{V"�Ió�\l"w�g|������BVb͸��Z\��7�ω�br�s�:�%<P����r��:@���\�T~�	0�0p7��>�~�*&&�k�d���ڠ��R\��a|�*��#mW�]��c�_6�6�ҏ�ޝkc���g�ƞ<���WGӂ�<Z��#�/y��PR��t$SԢ��*�X@bo��y}�y�A�f�{Ƭ���G�A�@��ɞ����oD���٘�
JZʥ��G�z �1K��@�	�u�~
�Lz
u�����fp��w��يIbL����DB�(�wt�Bw��o�>�/�#*��=�5	�J�1i�T��6}1�U�R�4���
�5/�4�u�(�;wW���/R�7��e����G�O� J����t��ZV���w͉p���5)g��_
�M�m���b{���3ʓ2J�����������}��ܚ��R�e\���AD��$�m���i�h\�]���Y����e(b¡�?Z�dh���r����G`ZD6�E�$���c��E����7��n�@��:qb����o|�_g�0�:��#���{�[-�&�+�j��Gg����Q�?�4�Y5�x����� ko����]�_��������6 FVy����,U'07\%\?4놗��T<�W�3��/2	nG�:��C�>}.����w���q� /�$?G����]x�<,#�tt�"�������EE��{�<�����	�
	bE�����^2�����/'�[f&6Q���kw�v�����_4��_�~�1�U�L�3Z*7�3�4$ѻ�iX���'��3`��𻫒���d��Zl��^�Iq�oݷ����i�= ��!.+�>�g�was��yK��Aֲ/b�ax��	qNv�e6�TYd�?@�5�M/aѺ�v����9��玙���-eiᡣ'"���X:�Z;W�����o��ټp���gS����o7����j��_�7���Ys�W��tF�mB�����j���t��}GA{��ǚ��#XV4"��n[Հl��4�k��]��_[Yˠ�|Sێ�*����p��@tC���u-�"؍��*� �d��Fj_ퟑ��`�=��bW�A*�)fU��Q�)���2{T\
�:lR_� ,���j~��P�?r��q:12�y5����)���=��w{x�l��aBW$]��L�KB�/\�Jw�޺�A!`�hn�5J�iaK 2pϕ���y��B���[����̉<읡�E�k�I���a��.�5ˬzp��y�-��dt��p�Z � ��?}B�궔��S�wQ����� /"O%�����@�r6,�Q@-���m-j��iu�]��-@h�N�m��d8�Ӹ����[���2(���#+ B��`�%��S�����$3����+y��&��(x���.���,��狱�#�039��5w�����%��������ɭk=��V5f��lIy
0ȷl�DT򩷼�pEe���E l���7\���_��u�[(�<7�K������������xC;D���x��/0����T�V��s?l�eT��Z$��)���:�Ƅ>���=��f�Z,s]�y|�]��mB0ƨ��i���y�e��\.���9{�e���{�պ��x�S+��h�pM`g��:��J|-��e�y
�Wt;O�*ꁻ�[�����!hp��^R�I��KL^v�STU�ʹ�xϯq�c��T�=�o��}�Uk�BW��{Кܗ���eu��u��4��B����go��$���8�2`ͮ�{��]k��rYo� �4�uc�B��Fz���d��M|���st�,�4���WI汓:�)Trɋ<k�e1�ڰN����d������pw���7�H�{�|D*��R	f��ܣ]�J/��}m)��Ө�]?>�1��J�l���y�&ߌ8Hdz�(�Z�ݏ
P��[?f!��)������@m�Ρ*��	w5H;��b�,~f��	�o:���N�sY��pQ
ʃ��A�
��X��h��1Ɂ��Eb2Yl�ǲ8����ɵ��X���:�ЮS�Q��,>���Q�J�E��[w��b��qfnXOvo��?=נt� ��%�o�G*�<g�`��۴? ��8&5��A,������Tg�nG��ٛ�L� ���)VN��ଈF����5�%06@��޾�P����!��W��)<�(KLJ[ :�1�X� -#AO�ģ@�c��E�/�b{Dh���/�{�VOQ�pڦE� hf"h�!�/Ah�=t����$�� Ǌ�*��L�`�S��!�E�\�F�
��N&����)Y"/�P�qD��j���<N	�k��8��$%�y�L]�r��3>�Zw��52K<jv����OCٰ���Vz5"�e�Aa���R�TS���1��@X.t���`�S�8�c��Bp�NA{sG�:���g�DjG���RZ�_p��F��N����� D`��-��2s>;P��G�iW�+7�}FAxa�t`���Nl�]��FZfY#8N�|�y�+�<8��I�+�1����%��V�.����C,fM��y��o޺3Z���H��^p6��$,��UALQo-}�4W)-3��o�H��h��dq���Y���g�	�i�Ҹ���Eq����|O6�lw�q�����H	�о��?�3�k3z���w"-
\3^ٻ]]?�s`�ąT�h�O2���� ���TO�T�a������@(3
~�o�=�n�ט(c�Y4�Q��঒�>�զ=��U�ʌ-�37oN��te�&g"�(6S�<��K��fS[�ٟI9_D%�����K�H&�!ef�N�]4��j�H.9a��Om�-���c�Yl �b�0��ϊ��w��D�����r�(bR!+�&�ҿ�@�NTA�t6߶�!nu��pu�Nۉ�MI$����?X�,�g��"(z!� ~�*���sC
8������X�W��xj��I��V�՞o8hx,ռ��]e^���Wi��.��Q�����y�l-fgiTFB�����mS�8&TR��a�Ȯ�$n3Uľ7t���ti�,|��2��;��s�#���8?O�c�ix�S*��N��N�5��4���-<ƥ�?�&23Y�r�̯�+_#�'�,O(E=hj�L-��?c������sv��p�����?Dyы�z,�+���$t^����e��{�?�y��}����߮7:��O�k{H���C�
&E���j���/�B�z����YR�M㈊�6v~dYI�t�Dm^�3�bW���i7*QL�.�����������	^��6)7�љf�+[���P���wLٷ�{n�~]�8�7j��]ʷe����a��V�b��M<�;�c$�8Q�􏈈q���~�&�d�p� ��%ࠩx�H���U�̉�!جZ�\C׋ǒ��IZPv֦�u���|�����_O�@d	�|=����R SdTpb�^Jyi�ҵ�tfu&O����f*��!�:� ��D�+�#۟;Oh�τm3�����R �zn3v�AYq^Yr�|�����F)��v�_4�蝒k���m�Xo�ʏ�xV:/����I�E,����^�wH�Dw}t���x3�ljje����>��3	UsW����*������쏜Z�K�f�Tl�F��z^��Ldp�1��TU���í3ۑ]���]}�Z7��HEN�j1f��h�V�`���D��Xm.��3���y/K7�	��q4�ֳ#��,�|1Sah>O�.j�k$<K�+ʷɏd{Ws���l���y2\��T�2�.JS�B�HaVU�c$�����@��C�jQXm�
����U��}zÐ�;��7.i��է����"����y)�}�c�NSk�s>t�`V k�o����oU���J �
m�C@��%Y�X�����A�R��$K]���
�*�bW�q�
=z�@#wIQqG&��г�I�s>|pvET�4��w�s�)����+�a���7�1?"�1��_<�L�M@�:�@�.������K�,��+L>L��T�>�u��j��Zi2���`G����?�ץ�X͌�PWI�X5/�j�/J��(ij>�u�T?�R��ֿ���m�ň�kerY)Q�P��B��83
����J,(Z2�Áv��E�]xh%�1%q����D̑��8�w&�X0������"���ʠh�"�Y�h:�(�4���hK���ޜ�<��	,5��3�豮ԟ�ܟ�{��o��O/��c�IZ��QzF(#�h��$O��8aݾ_�K7 �<����P�@�������]I�� ���ɑp5Е��z�.�j�e�S%%�N(N~E���^=n�$�/
Β#:��+y��QwX.�^��1\6�x,9G{.��p1���Gb�@k��wZ��tj�u�{sR0O����K]mW�wd��,�Hיb�Bk,m���}fE���D�mPy���b�bSgw۫�c_S>U��_��A�pvq�$�:����Q�+�����y��=g�����ƀ�|n<afB�ম��Q,UpU٠f!_>ڹ'�ii����#ּ�1����}�:1gT1
��m��ѿ�N�-r9�pF�l\G�툶���U-��9EEp�֒����Y��v��c6Y<^�F�/�"Sq��}�6�`��re��M�[$����r���QO Q �9�J���-kl��fp�a�0RhK0,/kE�j�\�:��A�Z�����烈M�7u��{�O�+�J��ilÇ-���*:T:��o2=O.|�����Vm���Ip�[KoAY�xQ%��"G��!`e��ѷ��Ӓ�q�j(�8��r_J/ͼs�o����7νK��Q*i�X�� �Od��^�Tw�?("�X�VY�w�����'�Թ?q���tܠ�1~׉SV�O�!ڡ=���Rp�%ਙ������<�VQ����1�ȏ
���J>L+�E�_���0.?��@���,]J�C/�k�awJJ��hO!��ϑN�����~���������K~"m�x��k����<��8ʶo�p!/���R�KÓ%�2��"�֐�$fv�iu"����n�#[X�+�|R�}L~*T|��nڦ/��P	Y$1c����M?����,6?��I84�幄旯i��Z�5�B3:d'�����$z��U�CB��q/�>N"�޽� ��<�,�/A�S_i7KLޥ���8n+�D$����#H�K���A�#9hwpGI��E�9����	g����V�8V�)�P�d���v�h����൭d>���2_�`����$�v�mn�<l�4�xL�)Źe5��/^�� ��$��v�Y��o��lϪ��h�D�oJ��]�zh�T)
�kUp{��<���u�����&��J����#��,F`��H���>a2�Η����t�3��1st��$�Tn4�!��z�	�Q���+�3�,��W��>�/ �-�Z�D�6����rN��㈋�@w�5C�v���J�mMJ�?q5o���ɓ������Э4T8����b@��KŦ���j�;6]b6)9��UJ&�$6~���X~�	���+Z_K����6����T������ٮ4�������}�v�'/�-�O�b�B�v�j�&|��ˏ���3�{"��3�ô�bԬ����V�6v��׾�5I~���2��=64��<���7H�Vl=��՝/��|!�,�y7J�\�����I� ���TQ�i���(�FbP����`���(1�D;��6�O��a��$�<�&��{ڴ���������Z����0�C��w�U�<�0�J5'l��:���M���l{5�z�N�]eV�%�e��5��pb�)j���ov�嗽�,��J�D;V�@A^���<�3�O{cFu�kf\��@^��3����L4��	�1���C���>�E��ڑ�ȕ�&�{���Λ ۯ�R��ʳ��ޑO3����	˱�1���ث>�i�`�s/��_����I:jn�X'�&�Y<_eM�C6I�$�[��~.��Ź��s�����*�P9w
`�-�Xr�X� �P��%C~3��������wV\�U���Ƞ�n����}�/�G"�4P�i��I���ւdI}s�l�d�降B`"��!NFv��A�~{$�Ձ�C3��H%�
���CR��B:a�:��9�nM�������h��YEM{��w����F���P��ie,Z2ѡ1]��0��|�Z��"	Y�kdE˂��Q���,,���ĩ�>/�� �P߸��@g�<�xə�y��a ���u%~/ha��]��P�+H6�K�!ES�p�F{j�,q-C��4F��p���
������fA��r��'?n�����S����I����0�NN"�[X3;���^0��wu��r��0f&8�E:�~yr\
��R3L�� *a���v�4��3�a�����d���=�ܸ0,�pNK�=����9�	�:IZ����	���ΧV�G7΅�K	9v�#����۝��7l2%�2Q���T�y�S��zb�;�'`�q�>���%��$�Lz*��<k9��� 
'����̧cV�����y>fG|ěL�F�Q���u~nV,���Ժ_<A%n�������q���2�VӍ(Y݆'Q�vo��bw�Q����ѷ�K ��vXMc�R�����Q2�͝8�_�|����l���9�$e�6Bs�����4�pݓWۼԅ-����]6$��{C�gE���, ��==!��^.3+��f4��PK]�0T'k��H�礧����:�?�T��o�@h?W�9C}��~�"��5�d�������0�Ӵq�>�Ӓ��괖��r�.��|1�۪x͒5etL7ǧ���@�ڍG/?
�S�)@V*�����\��8| �VlL>���@��/5�{�3��0�=�n"��":a�q��
��W����+��D�_g����^M~L��0��c�8����*t�Ʒ ����ϱd��j�?�h�x�٨tS&,�`3�P�\�����b,q`����wP+��Od���T��%�a�#N�{E�҉見\~�b$6ȿ�<%�Z�]��(��2_�g��70a�gzZGہ�bA��'e�o����Ms��/XdG�5˳�]�����=����谖b �؁�ր_x|��, lk��6 z�ڿ����М��A5M���x0��6qɂ���oé'<雞S�.��eC��+q#P~�>f����s�ZpY�$�R>��}���ſ� ��cr���.(Zn��u}�g�K�X⛛�7G)���M�F�G �v7����2O����x�����v�5�L�	Jo7�K�����h����Ơ�Dי�)���rɢ�^2B��S�nà�޽�<O�����l�V��o�&>�H�V��*��{��#j�.I�����ʁoeU\�re���ܔϦ���B^�>�����~���}��o��-��z�YUo���>�3���A|���8_큘��U��T�a� ,�Ƃ�.\)"�Q���c�yxo��-������Vpfʋ�O�V��/5._R/@��6��,���;��=�^&FX�^�q�\z�*�d�\<W���P�Z�oo`�o�v�����^Y�^k���ٜ�b�����xd�
�/3$TOq$�4�$���o�,��Tk�\ G/��5��m͋��I
�K��V���8�lp4S��4α�l��Ȥe�Ee��)4
0D6i�Y�H�{�> L���H���]�o�xF�̹A�M������L�'T�0*�s��
dN�	�|w���a_C���K�k6��F�Ru'�{@�g��dè^'f�'2�>'���)�v��WL y���7  �x�yƍ?u����n���p�e��r޶�a��%� ǍDA�h�;��Z�3L����%1*-�7	J"]RS
v�8m��hydT1!*MS[��/R!u�#���NA]z+��4��t�$l
����'�r�� \���f)~R�Z�5I�zӢ��m�?���e���B(��Z
��h���e~�\�!��
$�)�9�y��.z��Ȑ�^W�dխ�w
Ң�3��B}Q�H�>��H8�%��{�����]į����`c/�I��l��ݖq��*�@f�8Gw@��;½�p=�s�I'��T]v�%f���^y/��R�.n�@/jgG)�?=��
�^iҚ���R^9�U���m��%J�#?���cU�k�4.�M�Oɀ���=�M�	��lO�5` �ޜ鰸�>)K�8�����.!���e���4O�jgh�/Z�m�;�*E���R*I}�k�5c (���0R�⓯x.�Z���c�b�{�(�W�f��ڞ�aek�L�P����YV��|�_S��w�j�H���B�L��s"!	��@<�7ϑc)p�Պd��5�Չ����/���9�T�d}�tw����M�=�n��hN���٤�|�l�� G�Hع�f(\h5�U�C�gf��H�HA�o��{C�:5;��E�9�^��H�B5w��]�4�N�d�Nք�2zm����ɘrH� ���'q�$<�Ȋ-�	�NN��G�QUz�e�xY2=,H7���"��j��CF��`9@��yK��q��]M*����ܜή����SAK3���-��u�x�(���W���t"�N�����D��դH'�|�.�d���כ��Q�>|X������5��b*&.P�p�M���0Eٝ�ѕ{ԩe���χ�Ef-YR�03��)Z�Pc�XfV���ٽg�2��l�|W�9���=�������f��F�'��=�9�Q_;Ӊ�} 7� SJ��-E+�"�𥅫��<�n{�h���7v����Z祺�	�����'��(ш
T�t����92����K׳��l
��5D�5U��4nD���;����`��p����-pE@�I�u	[�cX=[� �Z��T��]�Ε�d3�>�ǐi�_�r�I�*G��'E<Ԅ�l~�~�c����[�=S�}����� ����m�͖�Od�(̤�,�"���'����H�e�ޔ���iP��1o*5�t�Q�ű�? ��h]9����)&%b�-�8��y�N����.�s�[�HP�4���>�C�����>��3b���h�WįxXDvIR�L*$�x�<��Op�`qQ��xn�E�eW�r���w�8�y^�T�|��2X�wh�D�Z��F��9��.�K6��Ѫ5ķKA��I��l��d��c2Cυ����Lt�8E��\��"Ngi�]����z��M���h09�x�gZ���PO߳5f�fV�5���|N�ۈ��Ô��:
$�ģ��r7|-�m�@��ܴ�38�����lc�+V!�]̃�Oa�`!M���K�9dsT���7	�WsD-�A��KS�8��tȜ�K�a"�/�oG�仨�[�}�C$�Z-�������C���u0Աֳ��s��o;�{�B̳�D��W�VY{��#�h95�:�S��&���U��*�������裋ī\����c�z|����$
m�ȶr���k�ȑ[�U\�Ҳ���?+��0a�;�KsF��SU:՗�y����"t߹�K-j5A�X���Du �?��:m�3�� ��Rwn��r�0�Bb �f�<����,�cV,���uK�C�L�Z�G}k�z-\6S��**�,C ����M�S�?�`Ć�	�-����2� �F"��}�u���MKu{��?��c-���?�u�[�h�2����V~O��簟��Ϡod��D�]o��l2�"{�N�ԆYp=�;z3���S#������v����E�;���;�@��������q�/��wa��f����0!��@PR���y=��H˩_]X��◽w��m�D񧡲Ȕ����G�Sio��$"Y7�9��
���HY�ҷz�
-{8Bh�?��G(��ݾ�j%ư��j����<_2�݊���+R�h<�j�_�9ڄ���[��[%���'�O�^A�E��B�pK�P9���>@�����:�xrr�2���d�%��)`h�����l+Vo��%���>��u��A��7-6l�߶��~�rND�����0�E��#=������Ȥ-}l� Ù!�dm1cqt#=}q|)ӅO�&�1�*���a�X���g߭�i3��)i�=�ɬVy-Tw�౛�g� ���u)x�q5�+�%��x6n&�r'P�|�}���~s�O<�~��(q��T��o��͢s 0�'�f$�R'>���ho\=?���up+�Q[��G� ���n�\��X"a�s�G�җ'��z&�Z��Ȗ��n=�����,�Ǩ[�He(��|�i�/�Zt��n�$����Y�Ѵ���j��*�] `�S�'�����&���P�Q��6��bP��t*]���:3ZK��[��J�}�}�bQHYSg��B�9�\���^
���J!��b��(�^($�9����e��֢��oM4
 �g��Su�ݟ�j���g����y-��b�Dgqڌ�9��� �,^�j'�@�=�J��*b��v�|e!�M���:��GlϤ�A�.�)vG2���*>�)(�0F�Yx��N��tGt�&������%2D~M�1�v�VAT�U�:��+E���͗U12�A0�A�&�HD�Լėu�Q@aӐ�M3>�i��|Ҥ@zH��1��4G[l�p���#|�&?S��z�U�.�z7q�N��|ԧ�9��x p���	|R�|-h����ד�����<��'�_Zg�MÑ����J��i�֩Mu��K��x���%�ONlώܟX��õ*�(~Fq$��y������5i�s��F�-�az8��@�is�3�]�ؗ�aK���z���7�Bp�$|d�~���f���"T
uvR�[������I���ɱ��>,
��_%��\��{5�E�_�HWF]��q���}#��*�4�c8�N՝�o�-������ȱ��5�;0bD����_daS)�lP�љpՈ+� �`����~<h�)	�/��?�)j�"*$���㟋�86�}�~�ae,*�[O�ƁH�Q���5|��χ" j;l*�jT*"�Ϲ�yq�.$����p����G� ��e~Ǽ	�9sP��}�|����� ���z�!ُ�X��{@|{0հ\��j�0k��SD�?�c�Lĩ<�5 j�i��3����#MY/��#z���E�&A�8�M�S$)�z#�&��6�;�gt��Fծ���K�Y��a����k�=�k��^|��j� u����*�ħ宔ol�Q����:�ɜ�}���f<�����L<�E�Q,�;P�&��] ���%��^�p�/'��z�0*�E�K�B��)�O�6�W��Q���EGjDկd��&��O�K���٫hJ�u�������+<%Z6m�3��`o�VE}�$Q\��U�Ř���o�!Wt��2z�>| �b�����7��l�RU �L���d����p�L;��w�yE��E;0<$�r����Yk�/�[�5-�"E@x�{f14Pp@w=��{^k�P�����Wۡ������}J�)���"hYøg����k�����X&`C�w�7~"ۥw�I##�ry�������F��}�#|uS��;?d�}��?���q��Dyi:�>�]�zJ���{{���V����������)�{} �[�i��*�e	��9~��"�柷��1C$f��x+2���ՓVpm�DtC���� zD;n��ix��$~|��{Q_Mc��Ӫ�xb���tB=�M�u[\(�_G�c��s��ŧЁ)�=Lk���H8=F���qD("_a��r��{�WQ�	�g��{���Y�m<i�E�"�ȺZ��K��8���$U���6�:�*~ _�gɨ��0���dH�>wo휸�W���Ǿ<wl���R�fF��>F��Փ��=����� ���wL|D���|n1��֙�:&�,i�D~ُ����U-��CW(
��-�*���	�������ЎJ�$
�;ΐ"D��s�N��ٶ$6�<�Yc�<A��T�Bas�n>-j3��K@�d�N�I�11�\�h��,G����h-� �H?Ws?J/V���V��"j-��i� ����fE5�������F#�pI-!|�1����0�e?�pW��%f�`?=��Θ���v�د��������ڜ�]KB��1<�Q ��_}D&��*+	5�y��t^�����9�R�⌻�`��i��rS�����=���ڤ]�0�߳5)�O<��Әk�1e���M���L暋���+�,,�f����}��D�[���Zc33��Nd�}����.������R��<z�'B.�!��^��hrf�#�����Ty�L-a��"��!Y`һR�� �9�Sa�]�g�>%^�~	�ހ��ɳA�����1_:%�l?�&ݮС
�w�.{�G�^��.6|��Q��� T��'���EM�47ZQ8>a�u��-/����عZ��F/�Yt�RX�l�����6���x�a�F웂L(�7P��Ʌ��(�y�\xB�O$ T|�#�.F��{�h>z��]ɰ��Ł�Fҟ嵘:³�=`؋Dy[-F�Ϟ�����P紐c3�$<W�J��r��-6�{Xh�*���A�ς�T~��~��\� Hԙ��n�3�NJ�9�2Ie�'և��-`�@"��y��9���Q��"����%��I�\_�c�Oq��6�LI��٥��O7�
!��tS�[��j�Y
�TM�� m��ם	�ߩ)�J�o$��bo�*a\�H����h�0�d�\ ʯ�5xɭ|�-��MA�FCu�!Vʃ�cR�?�nu�Nw�W9����;�c�:���d�5�$�n�"�8��A��c�������$붰N���a1L{D  -~F����8P�m��f��9�aU�b^� �p���r������x�Ie�I�(��O.�y��ĵ@Bj��*�`@Z��C�uX��ɃPM�l+��,=�y��	I:̉�"��
w���C�����cV!��V���{�'{`i��15�t�����U�P]-�G��-{����sJ�&m��`��l���O����=�g�6�ܧ�,�8-'ֻQ�eF���/���=fiA���A���Փ�>�= ]����q�"2��jz�N�1 i���pK��Q7?�1�M�z�5'�|�#�|n�{'����� @i�����	��A�����j4���ѵ�7�����>��|���R����Ғ}=�8􎪦�G@*D���i+D���c���xV[��W�;�!����\�+��-?��%�(i��$����7�Gi��a
 �� /]��ͽ�j.BP�M�i��7O��c)�3��X�����B9�nĞ!aB�O�J�3��y���%��S�;Mх�H��|C!Ŧ�k�[Z���k���:�|L�HzdO+r�s]b�ISU1���V >�Iʯ��Ggab����t��An^��3V,���W�Ɗ:�]7�+m�e�qB0}���;�N��Y�c(Kd�^�V���v��D�?rkܕu��c�>����7����@\�s�%�JE�U�J��a�N�*�7�����q�P��ɨk͒t�/̎��l�����C���z�Ȟ�1 ��a�Eh(+i�������qO�����^d���Z�j�?���D�u'��w�Z���䏰�oZbAwoΓ 7�#�.�A=���SJ�AA>B�*#�|�G�ITQ�|��m�*)���(m8�H����"!��aA����Oa�Z����B�|H�0�o��u�Qm2H~��%x�Mz�
�QE�,ǯ��U���b����!���\\��G���@�W�Qj�$:��-~&yx6��V*i0��Qg��~E�7���ɤ�-x�(��׶�!�M��~��á�.xS��h��B�Q�S�,9�*�i���D}�� 0�?_%����@�YR�뢦�����>���
مzo�����BFgF��O]��B����3-������ۦdC(�.������0�6���o����
��Aw��ې���ָNE�h�^�Ӏ�Ο���r�0���
�8�����P�0b�6c�ƽa�y�h5��bG��b���O��*�"Dd���N����<֯�=�ӃgeG�)��<�����?�1@�=#m��B��}d��]�&��Z� T���3YF�fd[j�K���̈́�,��w��X=3*��(lZ�2��n�`r;����O�rK�I��C���� |�Χ��х���:��_|{!���6Y>�k�Z�dq[lf�a���W��c!��6"%3���A܁�ç��c+�%�l/*H1�cV�M�UT�M����pe�%^$g ��.��2��{�+���r��:����+�r��|͋dlF��G��Ǫ*�����6ɚҋ'����P�V�F���"_��C����C?ѱ���[�� ���"�LLآ�͚Bi�9��R������~����:�ܡ���:������Bz� ����<��ʋ�t�up�x�(�9���#d���$���*B{mh!�4�]��_~�s���:�-{���~��drv��"g�5�9���+ȑ�p���G�SHg�~ �q������T���D��N�&���{/��8ݲ�T�{��W���
��}��������8��zM����X����C�`xH��2T�H�%T�Q��p\����;cE|`Er�RI�����Q�ʷ��_i���o�4��%G[�e�zQ2�5�Ȗޛ3�|�AK
Xc�2KL[J�iq��c�yS՟�OaN;:Eg�h?���+M�|�^�P̂\���ւC�)�4{��^�78�^X�HG9�+j�W��Tz7�����f��/J��)BH#>L�y�������Y��/��q	�F^��3��W��L2-�_�������OX�'Zk������B:��@��g�R�̡��u��(iX�XٌQ��o࿒0EnjK�@��ͪȁw�qET6���g��I{��#��G��c656b�b���D(�mD^��a�����{�W@q����ls���d�&{Ls���!��.�s��)������/?��:?����40)����<P`䧏���#ݨ�L�)��|��?���ʏ�1 0rC죰z (/?��L���ߗ@b���<x3J�����;���4Ḫ�a/���s��T ���6��.���������%ͬ��������۰�@�2;K�5����ch�j�sMbP��7�~�7��;����?0���(3~�֌4��������PJ�Q��b�:��XC���V1�!�`�?&+w��>��F(�߆5��LT� �,�qW9֋�5����O.�Eq3�E�"1�S�%�E$?��;�_���e�8��q-H��ǣ���WI�w��!-Z�ȝ�tܦ�6��zexI��sA�ε�I,�3���ϟ�*��'=�"Jx�� �eų@;�q��v��}��M�P8���R��/�X n/r�݊�2Z��/h#v(̇x�;7���J��$ �u���v�ˏ8MO��?㥑5'抳�����w�P���h�z`�iB�m���^�{pͽ8�q��9�̕�*,�+�>c!�d��1a]�E��@�R��_i2ϲ��~�w8��_}:�P�OZ �6"S���.ry����`vuY�v���L�k�ϟ���}|nn�28¬�2b���8pj�>�Ph�D$���7R9V���!�Pow�$CEU����M+o�#�OZ�j�i8z!��%:t��������ﶤD�_��?aHI9�'~��75�m#�����IMn_.S0Փ>��"�BN�c�P��*r�+r�Ko���&��?)ԲJ��.nG�3���@�� H4v�D8�_8b��x$�a�=�p
\
����q�`�2��JS���0�\1��УC��m�,��3'�~۵44�-n����uB�KY���JpH�'V�ze��z��*�r�k�x.����m�4�s���V6�e�#�^+�`�e�E2�ׁF.ҙ�7r@%�}͙n�����1D�	��*k����ʉ�.�7H^��"E�n�7�مޡ������'�iz{O���}���s��zU��m��l�~Kc��i���o�g��$��Q�3��\�l:O�Z��r��Y%X%Mg�2g/��4���B D�a�ֶyӄ�-M���E����I�[�Ac'��G�(ےyɀ��W��֠qAQ�A7nؕ��Z�b`���e��� �xj�B�ٖ��|��_~��c`DUr�IE�$iQ5rD�c��[�$���8>� #���"������*���3"�W�b�/�UAM碨8�����w,zO/�o!�x~��ՠT����B��E��q�5��b��I��4N�������n���ɂb��}��Pq�2*�9�<�.����!�#��bS�p���p/Vo8'�d-�໧���k���ʵy����^L��t|�	])`!�k};كP�ҍ��\���`�&N!	�>q��e;��ڛ�^hY���Y�����q��q	���G��=��_
Ãb�f؅/p���Q�XY�B��N���`B;i��S2��\.q*4���@�ࢁ�ќ2a�*�@�^�F�����ښ�F�eԐ���p��f�����J%�1/������a���B[���P1���7�y�A|4���:y��"qC�sxA{�}�ro&D��U጗�79	�MUuRc���tl�������h;�)5���g��y�ɺ�"�?�y�U���L�"����r�~��}L�콶8�#7�W�F;F�c�.@B����&��8{���9L�:bB��)F�O!F�Y�\��	�N���gvv�O^֠$3J(h8��B#HԺy`�?̿��q�b{G��r8R/��,#�~�>/h
�&7�0���83x�%��Y0�G:L+z���߂b2���jZ�`�+�c�t�Kɷl�JŇM/��)���QG���Ģ@t���vݒi\Yo�MS������xw�Q%����������8Ev�@ �ΕT��b<� >��SB�I?�Q!�{�V���(���w{⭧G�կ3P5 O+�*��O�ȓ��4�Ȉ�+���e���DG�f�I9�oFz� u�Y��($��`�Щw��GaG�`�{��3ɛ��شGTK�8���	����%�V?�		h�5�,�|��>jEM&�SX �6/͚�@q��CY�]�!�~S��"1]6w�:�3�,ü;�-��=Ƶ�Ş��C�U�y��j�Ln��O}�ڿ�p4<@�b�)=�%+����1o#��z�^&WO���ѣ��)/�- ���y?�2��@w�G����ٷ�x0��S����g�]��b���6��2�7�Փ�S�@��z�]�r��	�ڄ�-~�� ���®�NEv4fh���a� a��O�З�q�p�vі�a�p�G�r�)5���p�o�Q�`��.������G��U M��%\�
y�P#P����3 g�E��U�:ͭ|�؀Hu@{9�u9u���X��*�rʄwR��K��9����s��� Mh��׺�7N����i�(i�O�8���g,�T�τ 0-�b�{d��U�}��3�/�Y����p���A�*���Ҿ�znH<)�N��=n�hq����S�_'c8���(=��mqh�-��_f�EX�U��w�7@��R$w���\x�t�,��&Th�ΓM[㡟��C��
��3�N�Ȯ_��ŖZ{΁��E��YL-߸��u|b��?߮}.|��v =���M5�0d!q��������:���Q��e2�/v��'�6A����^G�>�A���G��u�̃$����I}T���I�Fǝi�� \%��|��:����U#%c�l�":!�e�#J��6��z<|��,Bz��?W3�g��^�p���ͶEi��Y�LH4d��h����UFT�$��*U|6�^ϲ��k�kLt�C���y����<TF���W+n������v&�`�H�#�0b�TY����US��U%@I^�������a�GJ����f?��'�x�?W��J|��^Q���vd1�� up�:&��^����Yc��N�uV 6�W�̘Ha�P�U�|�1y]-+ꯐ��Wj)E|Vq_I���rT�l�G.E!O�0�����	V��;��:`��\o^����;�9����U)� �ī�̮�k�э��oIS�{ :���49���߲���lqEF�Pt7�.�K!_�
z����@g�g�؜�'����� �Q0���H|W��U`Yr*4��e~^wxwR�Z�����}^P�Bܨ���F��> %ʛW	Y�k���>6Xv�K��j��;�3�׽��'$�u�f�ES���a�"'jt /*�@,�p�2x�!�v��������²��$\{s�zIw��a;J�B�x��q�D n��Ĭ��CS�N��ZK�l�����Pz6�t����Z!��C���HXND��y���6�0Cఎ����L23��L�([	�/�ջJ�ε�}�*&�4��j�L�*l����1bεX�/c+H"ջ�P���(#q��g��K��.��U���M�J�R#G�b^�\�U<b�P��|k�\���X���F�QUS~�'�|�Dk"(�>���ot�j���$�k�n��gZC�Sb[�ż��&�$R"�=kќ�~e���;�ׂ!�%�J�|�8�9{߆�
�!��̑=\E�1*�pJ~"��3ڈ[CY��s�A5�jgǭU��XЅ�}f�%뫉���)�(�޹Q7BLfh���TA Y`;�k�<���~U���J�ʿ�ؚ�V���dܯ�Ș�.��L�'*�=ekT�J)5��k.��"=��^KҼ��a��'\.���
{��R�	q�8R�M&�]r��N������q�;�\3[B8������so���e������W��#OxgP��o����J�E�_���]:�D��!��l1��l���e��x��a)UfpO��W8Xh]��'�6���F��u���0���A@E�2���G^�R��=!w��K��[��WVC���a�a�e�2W$q�+�/��|��r6��b�Wwݜ�"�	��V�I��M$P�P���&3�H����˘�#"�s�ʓ�хh^�F�s5�z�OR�4ߗ,|avNh��lSi�q�#^����c:Knk��(h �N����&ْ�Ǎ��{���-ڪ�"�6�0���ǆ����ݨ���	§��P,�N�R1 N���;z\���������	��_E^��������/��a'lMB�i6|u�W#��6����a�o�̞�K�~�Lg���m6�&����Z첝���z�H�čln���n8�L��9�ư��3T|x�����1%�[.�{��p��'(�4�a�d!Z]�ޡ"$�PD�@�� g-8�=D��ָ�,U��2��̓9��u0�=Ï�?Xth�/��7�P��}�p�t�U��$ͽ���2��8�y�x���	��6��}w����:9 *z�vi��X��5sm\��2�� ؀�8(�WIÌw� %j�����(�D~M�˜:j�G[x���lͽ��5�aU��d��t��
�c��^��P�7�p�����v����6y�~a:���S�h�����1�sjuL!	.��a_��˺�[f����|����������8xȨ4&�(u�\*$�-��A�q�Uʖ6����3�h�a���+��hH�Ӂ#�<���	�����aױџhX���Ni�)��rc�?ټ�ϔ�zv��LJ�&�6��;�ʮ^�<����d*���>�"���p	�5�h���H[m�H�+�Z�N!�(�M�Z1�f���7V~4�����k4��_<E���}�d����D�r�Bi�"�~�n�d���n��,���.~������/��q�$`���:*/ݓ��KڢI��|,�`���|�n��R��:P��u� �V+���j�������e:��R��D�;o<��,d��'�,�;��w3�%Pd�9��k���e�wM�رQ]"�����3C��d�e�^L��2�b)��	��'R������3:�&�3\�J.�MFܒ�>�!��罝�N��Q�Q:8%�5k���|o�"�U����b�|�3��81�ɛ��t��<��mL�q�R�h�%pF�<U��ҵ�����$�'+>�rq�O!�0H]5+�L�*9�x�{2�q��5�ܭEeo`�S,��?���6�C�TW�`��X���C�ӸS�G�<�A�_�1�&��t*ѠVv��hF�}��Ʊ��9�1)2�_>_����m�`�����b�I����1���t�O^�����R�h�&!S!c8�zP�d����׽ ��Gn�j�N�%�f���kH�]$�k�Fy9�{*p^+�2�Щ��T���_s�N$%�n;�3>�������*%Z��骒�E��\U�x��!A���|,�%�:�X�&�4�ۆV{��c�y p@�gD`f�@�E�_�u߀��S������7�ls��
�i�k�^���ƾ���A�1O$t۞N�,ݙ{1y�^d�E���S"F���iB�����xH�,��:��;�}�[��T�3�Q�r���pj�(˵�tm9J-U���r���������m�bx�8}� ���6q��"��rb٬xE�l��R��~�C�tau�d2mF�v�d!����(W��ý\��y�N�������o׋&�w�8p�-x��)� �"���h�1oD�x61S\�;o9�b.ۣ;�� ���s��K�X�Ͱ^`��ɩ�̴wXB�=v��̦�
��~Tp:���A��$�DJ��ꯅv�
����q����m���BPoI䑣8p4��T�+��'�5��q7p�,��m��M�S��{&w,Cu��U5E�U��xH�h���q�ѓ}Q��.[m����_魣���|�=M`1�}�;����]����1p�ؿ⎰<*ϕY�X���}ʬ�-A��MZ������eW�O��GJ`�~u�)����1�Q�3&;����M��^]n{A#}��T��¿���mR��Qq})��GLN��0:	]W�O�q��*�����	��h,�9��p��4�.vE0徺�.��)/$ӆ�в��<b�/<(��u�����>��]�y��D-íJ�T��	�-g%���������6K�n�PyN�j��u��O(!4��S̹�V�!�wb�!]DxM��&nJN���V��<hu�[��>�6�qn��*�z�����N5���α~!(�@��z�h��`a@b���)7�[��/�����yF�)yn�I�f�k�����.�+�hz���Yɧwl��j�rP�"��ä�
��pJ=�g�WB�u���:�7�/�,&}xb?z�Mm��}6Hm����J��K�3ߗ�f� OV�eR�3WK��87[kz��J�]~m0o�����J�^hջ\�W�š{8��m)SZ���������g�!�����O��I\N�=r=�ʫ�Xߘ4�h��ܢ�9������P6|F\��q�JK�-v�Q��G�uwe3 @��h���v���0�~��jh�^�g�<S�R�#�ӫ�\u�����`�m�K��s�z?�-��@��&��Q�5��@����N�Õ���)��~1�f�	Y�z�HV���-��6�´������%��E6S�������� I�u#]Ņ������b(�ޱF�	���Z��0���*}V�}��ߨ�u^^�!�9M1
Ƣ5�=)W��Rg_����e��i�w�mĻ��q����}3 ���b��:�I����w@m���B=�m�%�MCvbvB\�a����̱�I�MH��8�����Ik�<x|�, �
_0?r�V��x@ks'���5�k��F�+0W�ac��QoE��l%�a���J_�q2�|���*mvY�ޣ�OwE�ë;y�A��i~qp-�֣A|�נ��m_�="�i-	GLo[��x��X$rg��#�3iX&�;���s��-���^�V�s�dZu��M톐��f`u�jf^��+���N?qg-hO]VU��G�)��<ab"�d��!k�6
�H糶�Jn2 �\Qj��[���2gZ���.7 9�^�w��9��{��{ͼ�A��Jx'0e����nV'�����y{z����Ny�`$��!r�.)3��b����i?�}E��=[�^y���Q������u�8���xn��:s/ͻɽ��g�b]�Ø�שٻ4k�Z=���h���)���)0� �OW��Z~��x#���[U��� ��8��ZZS��M��r���(��~8A���p}~<�ʿ�H9�eN��I�E�g��"��-LWj�ev��%j�_�ǟ@k&��	�X�L{R\���!�U�	�g�V�b�Gyh���-�*+O�m��)b7)�XX�k@�t!}�f�~�e�୴L�miM^56wģ�_o���Qj�!3��
6`п��΅�)�m:4��O�	{���d^� �������|ɻ���Ow;;\zd����t���I?��͎7�C�M���?�Ra:q0���D���k�e������=	ކ��r^�<k�d,��:������O�x���ĊH�o�b��.�@�5%;g���]���g$�uW��Mʃ.�+�h��RX6�X���QT�c���T̷� s��8���pB�>���p	pX������y�j��G���ה�j�}��zT���6HEj\>�dp�� �@�fŬ���e� m6,�O�aO5��������)u�i����.{?s�}�}^k��HNjo��@�l9�ǧu�(T�/4~ϤC��0Wr�~L���v�˺��(��:8�}5�
_��ڤsz�4R�Z�Րb}ip�#L��f�t}����,E:מ[��[毝h�H�p@�,�_LO�~X$^�[��M;*#�4�XہW�_�s<�]e`b[�ܶ)��EM�탍^�Ņ)f�W�0��� �w�ɹ'P@q(֕�*rr���{V?��ק^&�+�!�▖QB�r��QQ��	�I�p�߈3��|�e���O]�[�9/ɵy���2Ju�E��K�3�1�0)�oew"�t�4 ވ��[�.�CP���@M�RL��X��S��N'#����dsI�T�!2i���G(��+\,�&Ug�|m�#�	B��X%ҴL����o8��&/M�WH7f���_*�. ;��S<P�if>*�����>�b�P�i�|6��{�I[Y`]mN���p��ʝ����r:ʦ�Y�����aJ��#�]� �NBA�{�AҺ�2's�d��Ϳ{% Kp�Z����?F��-������s�X��P=g΢��U>� ��֗��^�ts�� ��>��Ƅ����T��J��>�,�j�G�ê	��*I���3*�V�zv
�U�X�vm����q3�(�e�zkܷڄ"ev��G����0O�+�t�$��?֯Tŭ�8�|�d!t͚��#>Q,<Y����}�Ǚ��f-^Yφ��g�����^s\�/""�D���+%df�]�$Fd��^4���<'o=�s|�i��f�(�+a�cf�hॠ�F�>����)��N��ǵn��)uk�0s�=z�;�8&}�KĠ��l4�S �K���L"(�C��*z�Q�}�9 ,<�I���z o=�v��o�8�'㩤a/{����HqG'I&���I��ʂ_���p��[��)�A���謓�AZ�*��Y@a�Nk2?9��̑�^vӤ��F�Ú�y
i/�<�
�"���<bJ�<]�q.�ܣ��[���1g�ͬԌ(�����]~ �q5ۃo|H�9l�č�8��s&�\,PKFI�]ŕ	$]�NrX��J�~�?���C���t,ļ��"�׀�+hf����mΰ������1�ȏ(An ��r$�� � 7v\�L-8�/����QD���D�i�v�Y���M�L�&b���1��u�+:�[^�WY��za�x�=��ֽ�ף=���Әx�9C6��i��b�?�f��F�զ0S<�?� �@��\�@|�̷�6�/��<�Aua��S�MF��o���!���s>��l����l��">O���|N�js_8:���;���,��[�P�ux�MlC�(��eN̙� R%�X����E]e��|�U�9t�l�!�V��+��<�C�! ��.rEx�4��(T�m\C�g�C,�4��#�+��|�������P�b7��"������"���ͳ\0ox��X^��G'(� ���wZc�����Ryc��_FV�y�mo6��ʥ@�Jfr�JJ�Z ��C�)"Z���w���<Ha7���e�䑾��������U��{6���r��6��-.�D��|�#2kEds�m�ߜK4�si�s��PJ)`Q�8ֶ�k�9>�MLεR/��Xr��z ��)��.��N��E[fܓh
��2�D��X�'����6�I�=j��ĀlD[�&��J�@z���h���&���jt��7R�p�N<�'����S�lW�d�Ѓ�PʬQȾ��207
��N�z?� ��g��ʧ�}p��P��"Puu�R���O�Z?G	@�J�h>����"<���2����n��:��5��!g���U�;���F9�v�� �G��D(���,Dtu��G�!Rs��8���+呙��^ߣ���I$~&�Y�7�
��ڙj(Phe
��m=��7Ѹ2����ޞk�q�-��O��W�@�AA�/�>�P�O��_����8�ŷ�޷�f�����^�f�OSW3�?�j����tR~	er��6i�������w2B���z�^���>04�oY�,c���\͉/��J�h���YT��f�����I?}�E���޻Ý�Q��Ӭ�Z<��� ���Qx1�)����G�<l���|�b�v��<+���e^(oT�2H���9��?l�#����z�<<m^4F�%}��P_�byZb�g#¦�J���)���}��a���'>�E
��E���[|���B����5�M�bD4�v*T���\���D�V�9�?g��,�Ux���fF����ː�QB
�+�7E:t�qPJ�B(�+y������
3E����� ���b�'����G_���CV���rR��%��}���M.���3��i���MU?�U�Ìx�Ll y%��Z3����5�*ܺAZ�Y��d�J-!�W+�{^^��3q�u�S�?e��鲞�	��ҴW��;�F�El��Y�K�pk��dVV3\�#v|�L�	Uǘ��ʎl,Cm=><�5�3mp���bY�^E.��0tY�&5��$	�1�)0z���)N���A�W��,D��l�#{6?J�.��J�X�^�Ȟ��?�������W��lo#�HKg��U�u��`L:��E�����Rw�1R�!dj)�%[	|�ڙ����gT��RtOzI�a^�Aꛨ٦��1�����e��p��!F�J>��;x�ҞL�<�MT���^rs_π{	��8 i����U�c@L��Dv��3Q��ô(��V�M���������{D�̬�Vr))�D�
P���̳�#��VG&3Q`��w7�����Ԩ(K�][-[�vBI�Q;��~$�׎5�3�����\�"��B�s�Ի!���/��[�C��s�B�Z���co������[#���7C$�Q.��fE5�_09V/�WM莰|��(��#�����<��-4�q��ֈ�V'��8�2�F��I\����&R򹝇�B�6�����k��U�S��>�j1V(M�9���J�Yb���\ *�%��Й�D�e��f��ה����̔z����Ż	G��8��%>A�hO�7`�J�e�?o\�v�H�Խ+��
F�9$y�=i'|��<0l�rz��en��Bp�6zV�@�p��v{�=�_ �5�&�D)��
�.w+��wM \��H��͢��=��ƾ$0[���
=����������W瀂;,��`��'z��h�K��P����W�8�e#J�y6��4	My�P�� dZ%���ҾK�跙4\
�m� �����7�W>6l�O�my�955J�IG���L�޹t�x���$CWZ���-�X��9A���b��b�]T��P$+/���r��X��_���^���H�rk�q����̢�r�?�z��z���Fj�x�����J��H����r���J1��h5*���Q�s8v��$^GD�"�D����i�9#�@ͽ����KL�N�!]�CV�T^9���;ʒN_�m]����Bj�i1v��:yD߅5�_|@q<@>b��6�4r;�}C�1����e�p0$����F�/�K��%�N{���������5����9��;�����oB�Ȼ��9��7m��J�����ɫ��_�ҥ��Y_�o�F�f@e�=3tF"��R���t#��{r�������4��|��Ԫ�;�B	F�v��V��>9�!�A"���>�迀Gp���҂`���p`���8��5�
�xMN��	O�]��f�ZU��AZ6�#�yI��X�{�M\,= (>^�����s�~n�NcH��o-��o�u�������hv3�s��SN���]x����Ce������Ԗ� �Z��k��|�CV2��a�!W-���Vo�"$��+�IW}2^�-0����NV�4���(y���0������(��L�'?��� P)�?#�����k�(M �-���
�@{���&�K�����@�_��3[�Hf 5�v�0Z������0���t�/��� M��� *e3Ef.m�˒���_;��^�Q1z~�G��m���+	���$�b��Q~���1]�g5���Mn�R�b|���:S�Ҫ�.D���6D�nĚ��b���z��Y�#��X{n�a�gl$h��w�&fx79,�������O2b���p�*�eT��U6x4?�[J������K��kJ�s;r��y%�H�s�l'��M��m��«aƭ����AI�i>S?�̮|�{��Pۺ��V��(��$�]c�E0+����]��t�Cm\r<\��+�vk���!�}q�_����6��yͮCT����C����d��"�s�����zX%��	V��A���~SO����I@��V^���dU_>\Om/�_���
?�ϒ�MR�{�}�_�I�r�?���)U����m���l�22���=;���h�P�={�����>j�KLO\э�(b^d>��q��{�,Q��/M?�ē�����/����y&L6�`��%����Ӏ]���(%�\��|���6���}��O�z=c���evh�9���-�>�[[�DLJ`O�=/;�A�
��M鍰	����)RU-Q�`.J�飃i@��bO�*���Y�J����M ��[Z�~+�� �j�J>�W�"qnYoح��-�KM��[�bށ�T�!n� �!g����̕�5e½�vS��A�U�*&ע�?4Iɐ�&x�:����DtPV��1�J�
.bG�X��� 'z�$�P��������%�M���p�ǭ-a�&��l�h�6��)y�?�نߍ�7�C�9�dch��F����������3��j�������BcU�,M��S�~���R�L~3�8X�̺�DR�A��︎[b�gccNel�ǖ�`������ɣ�O�~�n���l��@Zs�K�U��.�l��<��4��{�#�!G�g��6�Yk��"1���&�h�{`��&n�}:�*�/'j�������k���}Q�� S��Z%pR�o�Ow0c5�@~����S,C�l�O_"���~3:n��f(�bT)�G%� k�^��"t��`2���ln�Y���@E��W�������풷�����J���x,N�5���E�٤�����mO�>�����;MF�ʂ���B���J[���s\;�\-��zy
����)5g�?� �w��b)��!!�p���:�W�^�ȟ ����{��E!���Y�&lݶ���KD�U!'��R�=�Y�p�����N�X�`�.�(�WMg���2�gW!u����<о���f�z|�?��f�m���`YP���J���Q�fj�s�RȞTu�GU��`�Q60.B�<j{�e
ۦ�.]��!h��g�+�ƣ�%�MQ���a3���`�����ekz�8����8nâ�{��L�S��6�d=jZ���@�~��\����b��� ���c'��880VU��Uv�~b@7����PX��e�GzP}� ��0�;��(N�ٽ��i����0���D��J�
�SV]�q�4�Q�2���gc
�0��nڃW�N��筏�OS��p�/'t�JW鷀���yf�55gձ�N��x�;B����l�;z�e%� ���	ߦ&�" 7\��j5&���/�S۴��T@tF6��V�1-����yEK{8�0z����6���->j8B��+��<�ٰ�PT���w�*A��|�Ie>��C9�<Z.�px9���	+C�?�ά��p��?_��7�P$ �H[s{N�ԉw��x�_N�P_\\ uR��#q��~��� 	a�<�|.���NS(�̚/~m�M�l@�j#�m�8�u;���0�,v�F	m���f�.�!7��I�T���O�g~!L\��b.�;E�\�u�ztu��y�p��F'�
$��V��ow�5�σ��3x΂_5��ۅ�Ol��(�H�9T���I*��ND�@ ��h3�>+[N��!S��jZ�����Dj��L��^�����}\C�5��շ��	��u���MW���d��+݈�M�B�+�����ƞ�`�g��<�K��I�Y�N��q�:��"����,Yk=�jUV��Cpa�σk��z�w��@���*Z̖�I�YVЫeMn���j�\��3�R.pN���H�97bx��]?s12ۡϩ���h`P�bf-ؼQI[0�T�Vݛ`pw|��B��y�1?R��W�)>dW`���]ZN�c%���������+���z����IZNُR
�B{��Xo!I�C.���M>i_2U��́�S��"��'A]��RN4b�K�	�Q���v��BaV�u�| +��OvFc�W�y8�?�}�9����$V5���1��_�́8.��_�����'vN/7��[CoԒ����u\o��ɗ4�
��f2+��A�ZqvmiѱEǵ|ڧQ��V�^�۝?R��k��&�
eVO���+Ƙ�%ܭ�ɤ/RS�W���^6�h�c���}M�J���ק�o|�}^�%� nP~��Mp�<��;Y�<9��{��NJ��>��Ԙ�r��nV{�'����Ŗ&P
?E�S:�5�'8�����_�w�����Zp��b�#�:>�d�ڝii+t�x*�(�[h������y�,�T1[Y��"��hc�y� ��p��}��� {g�?�;YP����y!4�<�$,�ƖZ�Ѥ�U���j�	���)&ISә�;��2�~��Ʋ���݆��K=�����U�(`~Z��ڴ�%X#a���g:�40����WK@	؊ص�Z�@?��UG��� �M�<�m�x�_6G���I��Lqor�<O,}}-�'��;J~��M�Ẹ�|���/C��E�}�M����i�H��%ʓ�y���R%2�c!��V)���ٳ�9�0@�+�6ߖ���^��5T
�\qW<�^-�p��4��Z6|��?�F����P�]��]��{���i�%����k���\�Ű>��	rޣ���=�r�0�N��~a��+�S��5��"N��Ǚ/�jPI'L%��"Z��;Gu4u�fg��/�ϔ��T}����$2G���s��q�!�7�G�巸���7P�"�4�f�F0�|\�P����$+6pkҸ�6�FZ�vq�WPt-AE�?�����	n�����3�S��dZ�.���PҦX椃E�W��%����ؽ�L�Ll/�[OS�n��5(�f3�����ܛH�H�z���s��?S"D�1Ԅp�V���=1Vm�f���S�w�7�t����Dm,��,����-��Z�l݀%�:�i�ԃ \��c��s�@˟�Z��xY	U4~1��F�8hW�R�����~�]:� �*���]u�?��Cv.��s��_a�����08.`��b'O��m��2��=�##'��x<�AoP������tZ	��N�����C���E�n�\O�mſq����F�6*��t�<TU�E$h�?��a���:�O�xN��f�����6�i��:��7n�"o��b(�uP��m�X(��u�z�U�x�h4CL�_5q�D�)"[�#�#n���pm��˘�_�a4T>��қ��,5d�u�e��{/]��
���"�*c���2����=a�F�A�V��S�0ڬ%p����K���EISS�f
�(ٙ��şo,���ݰݍꠅ�����_��(����&�{ٔ�������7����R{��X�{d8g�ͭz�`;�Q� ��|��w����ܙx:�Y�	��l��f1�m�T]������m��Tb�oR�@�넗�KQ���
�ӡ�`�Pk蚞_�}�C�g�dr{\-&�n��u�z2�1����_Q�K��|%'��E�r�7���]��g��y1��n6��(�o{�I}�]�}A�'Le6�,g܃YS�k%m�p�?ίJ�����o�@?%ػ����f�hD\��c�~��D���-j��``�ބ�.U/� c`B����;;B��t{�t ��KqF)(�0:���`�9�+N��G��́_r�xm��%�O�Dy�+�dl���p��H�LC	GK�F�_�p	_�y��*��f.��R�7�/���PN9)������^�|e��m����fg�E��D�!����p^�˅`Z(J��}�{*�[x)>��(�i�ʡ�E��]؉TN:u?��?�{���&=`���S���:7=���k�N,����Z�x�a���}��$v�+�(S)�I�1�W�E��`F/�t��1�ZKy����O�6��R$ui�J!S��N��F@h������l��yd���b4c�*��z[o���?���
k;������8�)��=������^��8��Sp�z/�@Ff�S �:GW�QV��ɞ�>7�����V����(Vׇ�,�̭>�pS\���= )��Z�<:���ȑ՘#��M� ^%���m�=в��̈U�V=���ݹ!o���F��!
�b(ǚz�2�1,����H͛g�\ϱ�bK���.֖�<�i�e�6�A��ܵ���c���
�)�f���0�⌃j�riݢ�_;�T��/��jʮ�P	N�m�6�Eq����V'�#�nr_�7Ur���o0��݁������wb�q*�2�Y�@����"}ލ"�۬�Q5S��&?��v-SM��q�m-�_���r �_u�m ��/I#�����J�Gʅ"0$X������k ��Gg�[��k�4���r23�r�(��E�	Z9Y߲Hַ �$ ���⟊	 j̫ѩ �n���E=I=��1յ�m����+����g|h`-s���Ņ�"F�K������^@w�պ�  �5�a���x6XS2_(]Y��γ�L$��2)��Y -�����҇�r=��������mF��&_�$�7��;'=��rሄ7����A��0�hu<V�r~�u��z�7�Ź%GA�$c(�ߦ��p\���8�@�kYF��-L������S�����5�@���=������V�qޔd������ԹdaV���wY�̷]�]�й_jX���<T,�\���y=^����� �_���S"�*�oM��w�I0*+%-(?���f��cڷ���8�W6���)��֮#�J�]x*�o��_uDvR׮fT �Ъ(!컴X�opwm@DP�m��Q��ME���>���˪"d������U�I&ɑ�ܡ�����)-���p�"�@>�?�[N\Z鳟Vdq�@����ķ�A�d�jA0���~��46X��GJ�/BE&��P��(�G\�MA�7����|_�л���m[dtk�+OW���n�F;��KJ����W�o;O�qy�g L��)�\s�*C~j�: ��Xa0�x&(P��(��#b8��Sl`����36i�-�<��ػ�ԭW�SCe#�w^f�zE�;r�Dq50��3?(5၊�~�ι*�L���-`>�^?��ްU��<�R���sW��}�[B��XT���wQH����uЗ[��L�*�^*��a4u3@%"����o��S�[�1��������f��PZ.��
�8#l۠d���>��ͨ�+�DI�<�ab��Gި��@Mʞ�y�j�"�\�N�.a�#�=m�Z�Z�|o(6CC6���wcYX�{Vm��������L||gߙ��]��L�=��l��9��T�o 	��A�o1ci�������D[*�D?f%��� �ƅ�ط�$a�iM?�����W�;�͘�s�HFz�3O�ep��"{1��*�5����j8�M��ŏ����eݥ�
��*�Ȑ��[�˩a��:��/�(C/�IZ��T}��q�C��9�2�T�r'��gv��.��،�5��8¹���ٞ��o\۠�\MIx���N�`F�������"Y���?�;�5�Q=Ʃ�mTq:;�Ua��򀫡ʖ��;�#��g�Aሳ�Ta ��.�gŮ-�e����9�)EmA�yMa[��ֱ��!^�	�^�,v�k��ɭz��i��MyJ�]k+
Fb�4/D~�{��=zu/��]���?6���<f�C��)�
�-@���O����4_�1֯�ǍRQ�Us��PlY��,Ӻ}J�6.�\��+�yU@�ٜ���`�8�VU�}ϋ#O�޴.6�4�^�.�8v�݊f)�}?�=\�;dO���"����v���:��x��~֔�2�
@�~
���`�ɑ7�0\���K�Cxo�t����w2�A�pɻ��6������ۼ9)�#J�B�ov>ŋ�%�����z�;�.%$��s��}��Bs��I�ء� SX�$S�����t�S
�����R�8*��gx��g+�|.�J>�M
0	a��2�\�"L/J4x��&��C����HJXE�k��h��qX�n��+�I��C�����ωlc>�߈u�nI��N�6��VX/idi�f��oB- ��)�"�c=׳I}�m�����O��O��B}W�M�a�&W�yp�HA�-s)e��-�[�m�֓;�3
1�N�ث��ƈ�xYy��Z�W����\c8�|_���*4(�똼���s�
�R�qK���Y�#��7>Y�Y�~Q�n��L���b�S����nrĩc�׬{\8Y����u��$�I���;Q�-U�Ҵu8���"�Q޹4��1O1Tљ3�����nކēI��Q���!f��{S�O�x��l��$��5�l%�����E�XU�!'Q�Ϥ���kƏ��\�$H;�DS���藦�j'zc����2s��W�a��eA�5<�S�/�Ĕ���cd�5w�?�I.�Jqf����`�3�l>�eJ��0�u�q�D�,��ao�sݸm�"�����8�2��l����!ڏ88u���y��Dfi#-��S�4��ԾȘcm�N��0L��L7'e=�Ջ|snz�fJ�:�
}~H��'��n�V=�&�h���#[ʣ���A�uGt�_Y"k��e�.�O?��Q�����o1���j�[D�8TT�ʱ�qڢ�%F������_vS��B��C�d��+����=vm.��= ���>�����{|pw�{^�
Ջl��3)���]\iWƐ
݂Σ�~��_�)�f�R���z;�?_�����8��~���&)�F��]�X�b ڔ�5;�R�<)�����_ص�@哏�D��MU�P#�K�L��(�UM�	�j�g6NF([�l$L�%�1����Ոg�_ۺ:'���H�)j�D"UG���̸y&ߟ�oW�I��=�*a�	@R�J����"��(�X{��k�6�\ Q"B�6���Gi��ޮh��.��h:>��ۀG��1	v�W�_#�v���M��+�f�J�+`>��{�*g�kJx�j7mٮ4ze�����?9���^�[�[��>2%�E�l���P��F�(���U�_�(
�l1���LaZ`��M�����J���0N�k���;�f�f�ˡ�73�S�-�^q�n$ MibR2Mv���t2߫��N{�*#)$/��i�b����-S*��߳PH��\�֩�7O�r�-��"���7�?	�����J�`{��[�� hR�k͜!S�҃um�!�� 9�W�Wt����F�9/�%K�鵧O�N�9Ti"D�Ĵ �!�j�au�)nO`�EvOR��0�x�7=*� wRD�M�6k`�Ed�:�:����F^��d�x���L�*��tH�a*�ٚL.����)i�$���LK�!�}��e��j?K�RJ���p�����O�ꔲ6���/*�6�m��t�\��'4�+����\���#
Ē'�ޜﾏ��S�?��!&���g�>��1��Q<����5����q�3�f����Z�߃�<��zf��hp[]��գչ�}q�Fh@��4C ����Ϧ��b=�j^�]������Q�z�rv�SL�+V7�f��Ô���"6�n�)K��\Y\5�Q���+�ĭ'�� ��A�,7j�Z��/[J�Ԑj�e`���3U�Z]%t�1;C���i�1=�ٌ7�~4����S���P(Zoaa���%����0�����e]�!vǿ��"�s�%R�\)i�.q�4��t�9���F�E^i��Z��\���?VG����|��+UL^�>,Kztr*(^�N��0���'5얬G��	�2���"
s@��<=?��r��+�r�Iȃb�U��mÖ�"����bS��q\rS2�t��ר�� P�_�0N�ߥ5���y�S%�-�u�E����ޯ�Z&����4q]���/���Anɀ�2�#Kx`��h��	zm��PƑ��ӥ=>B����� ?
N���/��ug�۲��r*�+7�f����d�ͪb�*������-g-�ǉ>Ӟ� %8w:d�TJ�-��	�F�W�J<J"%��[}IJd��Saw��IҞ����P�-�,�j/�V�$���w�+K��H&v^��"���v[ֵG�t.���kl1ָ	�#�5��4��KG�%;�i�h�T��J��Vu=q�C]�_�~�����'e��i�)v�vq�˨�?
s_v�-f�t+�?���"g��#����ʥ �=J��z'��ߋ�b^�4�,�.f;��;���\7�*��$Բb�y�c~<����u�CtLJ�o���X����nlпL��ӗbЈ6��@�ͷ�2?R�����,{���(1x�V�*���?sa�U�oW��#߽K!�P0�\�@�f��XHګ��	o�f�����
��BB�@�<�����G��Ž����J��0�\�p-*�m`x��c�k�{>�&ru�0�'��������C�G��3)��uND�
��	���^�	�l9J[�e��z���u��C���g�zj ߆f=g�3�`�7���(���iX�^������F>�-��*�	m*8	S��C�ٞ�4jW[�� ��c�&q��	ϙ�k99�3�caMQ���=������C4�6�7#&��{�KPW>����顒�z��K��<�h��ǯ����E�dٗ�������%t�f�rK�Z!�4I��B������fu�'֧0|��M�Ǫ_�PjM����u����>YE)��>G�N�GR�c.���%���D��)҄��DU��Z�#lly u��1� ?�g����z���G �y�^���*z���� �5Iq?R"G����ͩ� \��83x�Y4&U���i:�ŏ�G����q��y�&��������R�?b�Ӆ#��dߢ�J��������m��zr�`z8dw� ЄC���2�w!��\��m�ޱ�� ��B�dƃU���]�F uve(7�Z�3G@q��4��sp��s�ӷp�A苐�?4�~�[gbQ���ގ��0���>k���n�[�f�g�G7�;~oH�xN� �O�Q- �:	@�M����]5*+g����ږ�|w�����ӬrOtĖjba��p!��N����c�,��f����T�\>!S��� n�%����#����B�㼬�E;��k��2&ϱ��n�3B/��7���Or�[��o�o���`�H�٥{�:,�U�ەI}�J>*��M�G�̻���4AZ���mڅ���5So�|��F�ġr3�hw�N�},؁����=řl`#������>A��>�����f�2�E�����X�y3���V�QD�9�ܴ��
ј�p��i����9��r*z�L�����g�(���b��]�u�����%�ga{��A�{��1 P���?���҅xc��e�?���
�=��c�G��s(mQG�i��0N0�!8���P"�bS���X<rhBa����H�wr�s�Z�Ã����Q>�E��ڐ���)2Aju��P�D?��&4?��O(۾460����g��܆�9��Dzv�=9g!����/�
�=�D��ϪiD�����������@:���ȸq�"�-�1O�]΂�=�f�%1� U�Ȟ�(I5�&c����d�O�+u�_ɏ���m��V5jf�h(Ą����$� ~t��>S�(��yD�=�᧍d���C"gcz3w������Eh2 ��Uy�	�S2]��=�8��- �]�c���7�����4ͫ�o{T+�&�_}x��]4�@/_T��SIT]�a?�y�W4I����|*�
&��T��a�2���j��t����hcoG.�d�n�lk-̀,�쌨e��!����W�p�H���Xƌ�9���o<ާ��I=���?O�b�y̠�#S)�C7WFf���D-1|X�o_��ƕ)�Pyw��W?_��X�懶���|�*��'R�sO����׵�08�k��I�|�t�����pU�!J���Ӈ7j�l�̖Y���82�	 �&��^�Ky{��Jm<4r��>5�V{�X}�����bh���xJAD.���9I-g� ��@����f����7⿳��	�Uox�cP�N���f#�D�CϱTM�&��-�h�Yr���2����f��pw�'��%oE�"�[ဂ��C	]\�z��Я��/�i���q��!��֏��ߙ�f�R-]mU��pȈ��JɊ��W��rP����5R\[OMՒ�K��O"�0Vs�L~�`}g���D��oT~���^F�n�����a��Z�4�v!��;Žjg�	w������I ��X?}Ay�R����f��#��mχk�~��x-'��1���d��9���P��xj)6�UG��1\�Y%{��qA�"2��%�<Opi��ޔ�,�~�
c��r8�L��E��&
�D��*$��S��8��?����(˽Du�礧���yy����TG<}
p�~��#M�[��ᒥ#X�A�
V��>G�����:x��_��

�U���&q="�����nȬ�}�f'�3-) ����u���7l��_}�J�c�I�\��Ե�OA<����Z��`�,m�f�	�1�BNp�<�BaJ��fD���`+%����x\�ˤ���&�U�����s����;�?�/�{��3�r�
�g~.�z1y�n�qsCh\@��O}.������zzϗQuyR̐6�͹�iƪhrt���R�RKEq1�*w��F�n�v��\��O~n�ݲ�H������M��Z�ǌ4Z�|���M6���@t�I�W{��2F%)��Il6d
��Yi���q�)U�1;��D���V)B�`<֗�A �O�-@��h���c�˴��}Dlo�ŢSKcZ�����gW�s�Κ���^B��"fK���.�d�O�2[����zN��8�s��M� ��x�� #�����~Μ)�N0q��W��2�dx۔�8�=1�+��7!ѝA\��˂��c�J��|�I$�L�o��{�FMƸ�I���-�Mw��8�25ø��a���P����n-R�&�;勉s��
��)p�*���������^$s���˨Or��7��}�AsK�X;^���Ë���VMlgT�U�7{?�)#�&���Πq��%|��.KUb� ��l��!c��<����E'~�����&��n��x��_�I�0I�Ro#�Y�7m��XYu�T�R���d���\�u��d�Z���x��D-���ý�L���lNh��/�����?m�Y,���o"K*�<���y_��ǽ�?�mu��L��
hG���h�d!}��ϒ ju�<�p��-S|��7�YP"�p��h��9��d�e�>�z^#zr�+m�x;��ՐD+���+r�lu��IaUȶ����5<q�,��aP��� �*�8���d1����&Uo�¬��h.�#�(N�O!���:.�3ޥ�te7��nt�,��l��g�oس���'����yZ��,�8�:6�v�ɡn�RǨ�|ޅ�3���E��q�O���
�LZ��u�Sb��dos�vH����V��Ȇw�;���O��r��Fx��m[4l���UM�\����!��X}�d>�ͬ�e=�\,k��{�?��_Ekb��-t�*���*���|��T�PgiDAo&�^�/9��B=HȞ6�9vТq��i����%T���j����f�rtu��`�֗ϯ�-Ȭ�X+$v�Z�nb+����f�9j�|��G^����Ǥ%O��git��Y |T:����_2�|�L��4��X��"+=��_³ Y/,}]�R5�ZQ�|§�Y� ����dnC�_�@o%��5S�],x+7;�]�(������5nإ�#jK[{:\���Fx�wǤ����g<��Nr:�]�e�q�(����>��tXS}r*HTEzi�)}�ro��"o�L����J�;��n��LmVԄ?����� �d|fn�0�B=���飥�Z���tu��u.@�C�x'��,$��x�Nt"�� �ՁV��UА�e񷲜�Q�C(L[Uk�Հ	�Y/�r8��X)������5��ĴO��iEq���9�|��x9CI;���o� ��.��$(����!����$r�C� 7f"Ыk�::ҺV�#����o����ƪ��Yݯ`����4��Û/^i6��[�St�}����*��oU��f��An�֧f�wIS��M�(M}:3��#�B>q�mQ'���$�����L��wx-�"�A�bo#��ԁaN��'+���O��a���T������t�,ߴԻ(��E��Q5L�V�oC
z����n�2���W��PpX�%���Vy�x��E�+��M���wA� �9���+�]i �<�W�,3�y|d]en�g��ٵk�'��j��܇.�3m����� �LC�"�Sc<m��3p�t���`�z���5F� ����F�K�x��C�N�_0�t<*�|�Oo�X,p2��kp����w�\�����P�[�u1�#�A[z��|$*���;ӌAq���Ӡ�u���-/���B�]7�VՐU)��a��Gd�@����/�P�a֞k��oɰfe��Nh��Y�C���8�����,+����g�?q�K�@BX�6��."M�ɲ}�9�]X��؛T�2��dP�k:8�/�c
�4�د_�b���?,/Á3��*!U�_̢�cR.�+r^z�aMq�)i7�����%-�E��Mr��,�.2Kg���6����	5���aqM�o��0��_����SH��t��L�\g'�ڙ��Ȍ�_����Ӷ#fjqL��]R3�o�t�T�x�x�T��pGAݴ������ C�@�)�2u�c��r[Bf5㶼O4��VG��RӨݩ����,x�=�Y�ɉ�H��V4s�,Hw|�j&�0w+g� *`D�1���	������N�g@
�D��Ы�e�3��.�7d"�z<�/Ý!�k��BN�ηʠlu�\�̘�=�������.���/�6Wjor�H�-�I¡�����������܃`e�C�g\�v��>a�Y#U'V�+Z�w&�y2��m��Q|�B��#��dz��*�߰�~��8���(�G���w��#��l?�a����h�;��!�{���Ro��&D��e����Wރ� �і${S���6H��9R��8ִ��%�ښǪ�D(�"�vߟ�ۥ��w�J:z������M�64��e���i2� �a�rx�W��E	��6xc�������N70� %��e�&���5_O�0c�ynG���?^-"-�x�4Bx�w2M�x���>�-IB�5�wU@�-q�+Jfl��q���4��j��!b)����v�'�
��Jv�c�}��<���xq���MLhy�hWh�v��w`P�v�|-?�rb���I�C�˷�����ZD�X�Ğ�;0L��4}I��v�])<���
�۵c��H�Ux�x ?�z�Y��X	k��K:�N��)�V�x��o���L�ٿ=����v�Lp�d�gk��e�*�GW0T��a��m�,�4��Cd��e^ �Csf�5�1�%��0��|���]��}���`Ij;�>R{q8U�E�L�X,SF���Z�n|���ʹjt]�m`�3{T���Vg��Y�h�+)e�\@qj���,C��M��o8��K�0�h74��>Ĥ��!��?0~������Vʸ�B�$s�KZp�<�:i% W�I#>����F2�{�`'[>#{( �/阽�e{���G!�`�d�0ً/��ݵq�!�.<�H���՝�5��g�{��;[�#;�D};��O��Z̢  d�B���̏=���Vy7�ҕ��DsC�a�|?��Ja�h� ��&]�D�=��#s��y_�������I���TX���00�(�0r���4ߛ�~{�(�|�;.���ns�U�(��J>�F^����]*�Y��� �{A��o��7���ti7q�Μm!	��/�z�LJ(��< �} �\1�$�1}��/�XH����e�x%n=��0�E���x;�bY�̪c&j�QVyw{���-30ʟn�}�9bz;�:Vi�B U��h�P�]�\R-~Q�%�Z_�c���*6ob������Uqk�w/S�$VP@��/���?�\���i����~��������7��M0��h���=�>���b���{�MM���PMJ~�(�~�E��*���B�:����H�gc���Z�g�����`�ظ��̙F�A�F[k$4��v:\�6*�ª��<f=�������5�6�n6U��{6��qq��l� �F���؉��"tpIq���q|y?Xw�2��q�Iw�����+�ES ��zmd
RO;Or�d�:���x^�x	!�c:줂�<��EgZ���u�2
�U�=�x������^���vw��A�+*�P!���;�C��4��Д1BB�a����|��<�'�X�ˋ�S@�AZ	E�������]ƛ����u��%6���r)���(^JyyQP�.��'P�b珸��׳6*a�������V�j�o���2iQ��u��N�R��} �ତB.K� ��$���V�ճO"�������$`����7�`ߛ��4���%���(�+l £<��
��y���RsKv���'
�w�����u�Ip~p��{l�бI�ȋ	%�b&?E���  bb�uJg������N�r�0��L��mm�J����]TGj	<Z9=l�n�6�rpd�q���L��3�6��+�9q��/�������ߩ쎪ڄss���&�U�\h �>��������yq��p~ϔg۰��c�RV@_L�f��e+��Sʣ��k0�;S:�]�B�T�[,�4*)�b���#BX���kU3H�z-�B�Jb��,�E%|�y�]�C��+-߃V]���--���>3'�� R�`x4��m��Տ^������Y�濋�-�j3�# �Ϭnپb�����)J�����+�WJ�*����ఄ9��2���J#H�gc��Y�����;Ω��I�B�J9��<�>�-��Z���N���ew��}Z�G�Ҋ��o�h�\̭jr�f@�J���b�df����D3�ݚ�a��q`�P�g�S0F� �Ї�q��o=�fG�_�S�{Y'SFr��^��b_�bC�bT���l�St����(c`�8R�Q����_���4J���rZ����k�#zAy~�v �G�y���!��)�i˸�׾�ڠ�R��W�������=��h����1Q&^���q#�#�#�ԯd-�د+�+b B��l�����ʹv�[~ω�Iq��)�c8:QB���4��!��̓��>G����M�X&I���X���#��#�������)����4�A�
�,�(�~5x�.��ݖ-i��GG�����і^S��i������齡4L���Bӵbؒ�o�W��FiF�0OwDX�2���\+g�'�� �sf������)��2�V+�
���r`V�/<��L�|�W�Td- `�ڝ�@����Ky_􄻱5��jM \}V�� =���P�-�z�$���/|i�{��6��y�%P�'����٤Gl�eC���H&� ����XE��P��/;��ח�x����%&T)��V�c>i'�Yw��I��\��v��S\���چ|b<�v������fmVFs����K�w��-?o�<�V���w����;���6��̫Ӏ�Ep!`E}����\��|1�qs��}�3%�����گ��;�r��2�����d�F��v%;Q���F��L~�'BMe��:���\����.q$֕Q��
�^]�5o"kk���n\�� _�;UrRP.¯�S���O
�!�?̰�zv˼g^����Ʊ��%�q�U�s$MЕ����_ϵ�%��9�y_���7�j&��h��XT���jy
-�0Oj�<t@�9����mg�AP���#)�e)Z���n� Ou��+W$K�o΢�o��f�O5@��¿�@ec�J
��sz�V2�\\y��o 0�p�	��8v"C���Ԡh�+$(�)w���[��*d3������<uH���H���AI�OG��*Uk��!�t�OPN,tyu�@"B�2�ڄc�X��7ݙ�����b�t^d��e����->C�²���e�|�Q�~�R�z�/l�饬O��OG�� 6�W��/o��E�_��"�K�Ǻ���������e��T��`Ձ��
v��7e�u���5u>��~���1�_ܾ:.o���7vD.���m��O��T���dl����դ��M{R�i��CI�����I�A�)O���[�و�P�.�T�;�1͑�ձ��=��uO��[C��̆��'�����^O�2+j�i�\f:�����J��x/��:��L��J�{��Y�-��m;��uS�?(��G:m�-!C����$�N׶H~�z��8�������]J�����b�;4V�K$K	�-��o�J�(9�� �Ly8{<}�O~ɩu�MQԛ�p���*�Ÿ�^ڵV ��g b�~��"���W���~}��]'
$��RJ�h���5��n���<M���㉵ ؓ"G8}�b�s��`%��ƿ}-�ofl��F�7��y�Kae�ȷmcݖ7�V�%/� �� ��k6?���0j�"�gijM�_��(�� �&�����J�e��B�Nu�Ay4vu���:�(I�S��Rx�/*#\�1�U��45�Q�β��r��IWu�!4�nЂp\�q��nS�鰸�0!/��UVc���D���ru�����E�̊�@������8!�Pr8�l�=����S/�|�\��j�r���d>u/���6)+GJ� )�����X�"��OX���oJ�,�̉K��t�}қ��m%��>�V3o���&)=ʶh%]N6�݆Me���eg�F4uEd׉�HBi� DF�y�Ė1eU@������q)���^�tk<4���3֛믔�u7ݾ9��������$~Cg��n���	L�!ԭU���-0�N 7i<c�|2b:]�n6`?��k����P��d���jU�A�!�t_ߋ�ҩJ~I�m���g�7���!n:�jZsØ�?��*�e��}�O�:����%V�wXz���o�23�嚣
h��1�S s��=X)�(��'�6�p^kv����J��p`���gl�]��A�l�'�׆:B��0��O��h�8��%~z`R�ϻN���7�]&���V*_���-p
�S�2��I��_�n�̈́f�nN��
���D�ֲ۟�&��:c�|�8��D�����o���w�)��{�i{]��n�q��?�GzI�S�����ْ̲"c�j��B� �
`���S4	d����Es=r�7}6f���:&�o� Kg�gD��F5�g���-�Xv�[�^Rh��� 1�8��Un� ��?	�`i� ��fތ�d�b?�Ä��d�qE�#O��*e6  5&���_�`a�\�`@vn�z�Hˣ����nQ�ɵ�5�FVxkB����\~5�����	H�U}��qӻ�P�?����!�!NE��-�����n���%\�35������sjr�״�1���Cj�펿n-
3qq�����;�8hZw@��3\��GZ�;gw����@ �J�$shy�� @4�OFs�{��o�6�q�a���������<DZ���Y�>��_�#]��@��#��>D�*WF�b$��?���W~�rR�p���}�x���_,
8��9�m]��a}r�;M��g�'�Hn�`i =�2KM�'�=�	���zV�	s�� ���-%�#`>.��ib��h�e��f�G_��5	p�lx?*V?��y��#O�����&�e�H�j2��0.�.�7�p�p�#{�������� H��M /ppp��X���D]��u�S�L>N���-�`u��4�ڿ&r��
^���/ۮ�.���o�C�|��ײkuuO�,ȶ�jٗ��Ue�>����Kq�E�-�*��{3}j���g��F7��Si+���oڳ�8P��F�v�ɹIi�S�W���n
|��s:y��niNZ�CE5� .f����M��J5�=�2�&� YSfo/QN�o���4o�W��Θ�/ >>��9���t>h��(�A�j�/��f:��v��9���mد?.�#��[�GҚ�ۊI�/��0uB�~x����SF�2����po@�Ӆ�3�_���8`C�F�9������$IP�;�mG�B#�K#�G�O����X��;ZH����kƲ/<<u����,r#��䰠��� ~ղ�0�l^��Š���A5��/����u<������"U+R�Ś��UkK'��}�H��{+X���Pq\x<��F���3��텯�)V�X�BALaP6io�=�RD,��]�V;�n=��&�6�F��k��	���~��ؓ����w,�KL�~t��m��YV{��D^T��Y��@�O@��\��Ƽ�H�s+����]tk�ȑ�k4W�S�>�ݑ�n$8'#��i����kS�n�L|Ċe�З����G���ç�c�/��XYG�E�|�¬	��޾��_w��"�5��;[��F�$������R����
f/��'�9q	gܸ|�s�4"ϣ��i���m��h�ک~\������s[)�0??�)1�S�jd����n�eW.�3^i�h�F�{�v�a��6�Y���o.�X�<$^��ج1	nO�����Y{F�[Bh/#�_W?F�7���%�"=�W<��q'�?8��b�u1\M|�����1UZ'1$�ۨ�����z����zz�㺈Ȱ6�ӄm�Z��Ш(�_��K���m:�h[V���Ls��+er��X�K�$�|?�Y��@���_[��Pbѫ�
UCw�����],��Q���G��xz��e��_/�l���k0EVE�����Z]�U���N-C��.-o>��B�� �����xk���->�Z*FcB
@1����������3	��)d!@�}�n��W�E>�����4�u��n�g�G8-�C��@��[�o� Zm��nY`/� ���|2!�e�(�oT,Fc�!Z���_=˦�6���v����c�]i���N�K�����[?���MG2�/�:�ӭ�������.���u�u�m��p�k�`���0���]w,ג��b��q�9{�Н~w�]7P�k�)G�I֒�{����0�t/{WqiLߣ��whD�!���G�(v[a����L~�ޙ�]΅	���t�0�핋���<ĮJ{j��p`.���T��؜�p��f-&n�(�Ґ:8���%��!�)|7Ћ�T��V�#�@nf�;�bE�2��-�M&[�v��)���,��w���������h�S@��{*���β_�4�p�#D�d��Y�C?
MŠ5�Jʑ�dmI�$B��}}��>B>,�a�[C_��@��S^:�|��w&
�@԰i ��14y��|�7���(���-�e���xlA�ډ6Y��u� P��/��ʏ�k���	��뛖	2�/6���.���z�J��V#����Z _�� ��r���f��|w��DN����`�E�O>�3�,�M�MB|p_�����SЈ�a���:!�	�^h���iᒑ�$�#�o�{1��j������W���a�P~�3�>AU3mƐ|�φ�^0!3hW�bZ�{i�~�QYm��^絵�����Q���{p�ϵ3�ͽk]4�q��1���ڼ��Bx�J����ץ1R���m�j�]��𷇚r��t$z"�j�z5zc"��:_���;f� W�z�~4�m�l������9g�iI-�W�{K�����bN�/{�W@���:0����776�2�Sn���E�&f��r�����M4�
�H��B9^+W*���j�ժ�$.���ˏ��.��%�[�y(ې,c��&g�B1�GG�W.�d�P��a2]�`&u�!E� �k��+�"�����F��4
�`�L&�TD�4x��ndŊ�B!���e�gh�1/�#_4���� r�	ȥ_a<�Ǟ1K�(iB@�zJ�ir�n*�G2�؞V�^�Z�o���حd��R�>����q��!����QET���b:DE����E�5��+������<|�(�Ռ
Ļ}-�e���	i��~�}m��O�Ŀ3��U��Իhڋ��U�VG���L�N��K��tU�bs~%�񕏮�%���!��1��]%"��� ����#9p�٦g��w51�H�L�/�I��e�Z�����-`��༕�u�sgbMc���\):O�k��n�ȪؙP�.�����H#�_�+���?2���J������M�����WR��m�x� _)�P�w�I ,l.O^'K
���3�8��Js�r��	�u?�� ���*
&�$ߔެ��G��G�Z�E�]��e�ߣ����zs8��6;�A�u���Y(���}�ؒ����<��S߀�u�ۖc��$9D?'��u-n&�-��.�Ѕ`"�4��^ֲe�78������!�^�Q���OT�ST��1�]�h�w᫥��t�'Մ��xZ���84>�$�	��S[H�d��l���9#ɰ_`k�x�`�5NRP�f̐C�9tƕ��87��ߒ�V��|m�R�Xs,�f�c>f���f��+������nk�o�2/����z�����c�E��KA}p:�Ŷ�����M!(g�W�1����筢��.Dd�Ɀc�sr� ��!]Wܒ�j�jz�/���#�cϘ���I��&�0���[YBhG��Fc�$��}��VW���]8=�JӰS�rŬ�^�������8 }���d5Y��So�Fœ�E�p냃��'�����_�k�L�����^ڟ���?Yrm`�L��rA�������Tv�����c�SG6E�nPo�-1�����%����&����CV��Cw�'�U�sq|�P�z@�B{�r�\�~UUqn�x��-��
4�߭GwC&T�Е'�����8lh[��������T&8ZP�9@�j}vZN��0���4�ꊾ�����M�e?^_S\�����:�򩾢��­[�$S�">��{r6�{�AtMI�"�j�!� �"d��[�"9�J�j�=K. k�g�h(D��������v�Q)����t׺č"Z�!ݦaV"��<w�v�6���_�q���vu|���?w���^�vG��;1�FQ�r�׷:�
��amfB��
����aa~aiL��6crD ��6�8����U}�ę�R:ÚWˬ�q�4J�*�]Ȼ�5۟z;�E͵�8�5S���ys��ڄ	�E�Cj�4#Na��_�����\`OC�b��J�B_�N�Bx�PP�Kt�2�
��ZQ^��L��v����0��7���H/�6:�@�f0y/�q�Ymn�6Jo�ԩ0I��x���SF��q������?=DIM�~��)ڕ���6�'2���{u��@�{<W��_���k��\����\;�qxn���)I�������w�tٹ��q�(S�v��p��UY�?|'lpyY���a�B&ւ	��L���dY�[�+C)'˴!�&��&f������6�_uYo��ױ+k�-e1��N�R�hS^1'���ҷd*X��ra��!�ߌ+�{U|>����Çl蝁�~d�'G�Z��>��p��;�\^��!%Ti%N|l`�n�d{���w>�������T��!�*��Í��<��ЎQ2Ќ�����YÊe� ��XET�e��8�{$�#-�P)�t�;}h/�5�m��T�v=:��O:kR��(r#$�̗Z�60e����.����1��LB�}y�\�~ j�5��e�݊(�e���4U���=�~�%�����s���|���F>���#�����R�����9�5ᱳ[Ϟ4v��H�v�g2f���V����#�K�y:j/���Z���U ���AA��Wd�Y���I���D�$��؛�`L�Ӱ�x��և(C9�'��^ڟ�출䀘�9W.��	i���gF܎�0���K�m�C{�۝�^��I��Cڛu������ۿد<9ÿ}�NÍ�ǆ�����	*0?Aq�J6&�U�Pe��
@)�4���ك���Rל:XoOK��Q_OO�^���]��3'&�W4����[a�qj�E�VY$�-�+�$�{�U���C�[�<�$�@W���?q� ��=(�L`������ƈE�	�gV{�U��X-�!�����4��߳��ʷS�[�c^���S7�Zn�����~O��N^����o+
8��f2\q��Z0l��_M�V�&���,�Z�L^ug)�s	��c�UY_��[Qɓ�#�����84�7�0v��"N��[���ä�������A��(���7������y̂��<�cBY���>��� �}Qc�&1������=�r�"9��]P�`T�=ݘ��	j�%���j��z��43�7� �4�|�Ɇ	����DVw���c@�wC^��X����?V��(��\��[�[yPL:LO.j4����"��x�Mu��cnf:kω�q�3�،f�2���R�?1�=��-p���mD�tݫ��ĔN|�/�KCO�/��:7@M}�Q��W�h�;���H1�-'g����|z�NF�Y�jv����!֔��!wU�v#9rM���Z�(�q�ϯ9�.a�.���Y�ǆ��ĳ� ��Lߨ%�x��@��\��	�ɷ@'�)�t����R,s�)��G:��D���
)�Z�x�?IM���m����A@���(.S�j��������2�3���S#�EG}�d�呾���=�U:��-y��dGQ�h�T��4y,�8۔�UM�H� ����&��D����1��Hس>�I�j����#��/!�G����m#W�nw
�ͭ[��EVm����q�]�0�vT&5yO�/`�*��u�L�^ʲ�1
��L��6u���CX/g���3(ԯ�0����+��q�$]?ou1q��zY��6��9V�O�뤡
r��#3z���W I��6��B/l	)aA��%�xST�«I)�����h�1�|�&�A��H#������d��b`�M�5�<�J���|k}�¦��1q�=a���V��$�I�è������p`O2��'�*�+����(�H�3%�q�?�JB������a��	g��P!���.���s5���ڇ��l��ك����]�������G��)���� Qe����n��i�q�����E>�����L�R��xE��6�g�4/�M���~���x���8IkK�q�p�8�F�ԏ#��c_��k��w}|@{;m[�w�ęD�Ne�QNO��0n�6Xb��J�:���{���iU>VZ#�@IJJ؄�����iZ�(��R���ٲ�c�T��h3[��n(�ҫ�M��D��߹BJ4iD���K�q27���Q��?���4.���jPI�hl7�ĜƢ�,g��Z;n� tRu�0�"����I�lE��|�V���U ������gr�]�d���=q�����2!�5�OO�͋� �P���J��dYǛ�^T��k�����/��)S�J��	�~{��拞��4��'�\����e���b��R�e�A±f�݋|�I��!bP��R�O�%((8���׬�ln7X3�G�|,������3��� [˅' 1�A(��� �.�+ܪ�"���#�orJ�X��dnOY_�E>�dy5��G��)� �R�#��DpN�PvC�9�w��R�T?i��vdjs�Y�&�0u���m����(}���)H��� _���np�ø��ʊ����w˲�)2��7�46��n�O�Ѣ�W��DS�"m&:G�7� ��K��׍���n7�X.��0��E����	��S�{-jW�d�c����XD ڞ��S�D��cO!��l��Y�_λer�%�b$9��1	�{��3՚�� /��Zt�����A��>B;1��6�m΍�qog�x�<I�ny-�W �2n���n�XR��(�n�ϡFUo���͏$���qw�8.���7���HN�M���@��ر���ϟW� :��,VPy�N	���k���+hQ�$��!7�mG�{"�O�"�"�<���'�o����%!;A�������G\�����Xt�i�����zSH��,4�R
����ot�W�W[�`#jl�ǖB֎���^��Ϻw0a3�HI]���Q�'��_�jAtJ'��7��[9<;��3�����J�
�F����g��Ca��$���Q�𭸍�S͛���]�肻Oƞj�d�WMP#�@#
�rB*æ�������Q�i�c��U�5��\銎�Q�8����\��.����P[f�t%+�<�v ���x�D�$?u~\z�ܘt0��+���>���Nr��R�H���a�&r���"��Tq�}��C�sB���^�ܹ�X�o$MVt���n�5��9bM�+���ך�����'����k�;�`��>_���#���V;�DA��i�$)��X��cn�� �=�͵�w#�] �w���h疣��hX#�l�on���ڰkV��r�1TS=����������3C��!E��lo��+
V�92�Hf�`�:���)�L!$'�G�<�?�E��{�%D��^ KW�saO�V��AU�+�{�!pBt]J2�#���6��=mN}!�!Eƞ,V&]�ZN��v�yGE����LJ��B+j!MB�`�ފX���N�S�e��;����$���w�k�[w,�<o���N�/YN]y��U�~�Fs��M_y�[]J�,�0~��c�R�vr�'�IM�YU���>ӂ\�A�.}��_p�A��}�3�J?��b�P�����M�� ��DE ��wMh�� �JE��}Cpk������#�����}vu�lK�4*�#=� j�@�%�N�+����pq�~��A�����Po�>0.{;�;+T��#�ySU�X{t±yW�Έ����z�^;�����W�g&��m?����:�����@r�����<뫺K���@�~6��|���$lHjG���}Z�3=�豵�)Dg��gs�rDף��A��^����}�����z(8G�qTB���}��:�WqPM�d��_���>�T���:�`^��
(�&��x��5�F��*����k��Y/a��v�Q߾�K����4XN9a��7w*��L&+C�h˝���^qD� Q��~�9VĊ��i�`�������j.�sKf�HY�2 ��7��O�gSHA5���c��a���U��6�~(�9��lh(e6?�9��@ck�5�b��7��&N'�>�2Sٮ������t5籑�C�a5�=
��#<��$1�ƒi�7|�)�Q��H�񮿼/�Q�%�fڅ9H
��贤~Y�eA�@9���J/W��
c�X�������~��I֖��]�ث/
h�k�/��)�|��7H�}�0�J�����)����-,<�`O>��ӥ��h�h��}Ik��I���Y&6���b7��u�<���}۽X��1 ���]���gUV	Eˡ�Cy}�8�,����,5?�����<_{&K��%�T'�8U�oN�Q|7C~|>�lJ.�YV6n��� �5Y�7���@	]ez�d�9Y8r+^�%���'K&�
��Fe=�*.
�)$G��nO�����.b�����m���BO����P���{��U��/�K�ϛy�(O+ÒYq�CV�.�:�M��<!����V���}�AQ���@�"#p��Vٸ�����)����)�ú�v���;r���WG���~��ˠ�R_�DG)���I�fn��x�
0_.�(=C�Z+9��X�#�F^_��m	;��B�0^.0��԰�u�i	�ۿ��$�3���~k7���Q�"�灎0��P�|O�{�����T��<����B�e�"�����L{H?��Vn |~N����W}�E�_�Hw�Ŕ�7�:XWœ�:H���x��TP���Ec3���V֋�Z'q�Q�P��n6)?ZC&����l˟jP_e���Y�Ծ���#��4$�v���F�r;YE�?7I�n#è�S'G��_Z����j����@Qe�}���1�Z`�q�LY�OV�F�i�G��1U�qK�����焴��\�3�ͻ~dw��豶�/T'�M]k>�~�X̮�fQEV[Ǳ)A�_�|ㄸl�mT�,��puF7��9'	G�ƣŨ�
86)�N z��DP����A�	��0m"�"�����0����5z����R[��)��d�R���ݙHz��@��i���>6��C�[�`�J(I�?�}1!P��0��*9�z̿�x8�6��A���X�d�ޠ����A��'�S�E=���m��V�JW���4� ���W`Pohi�խX����3A�h9�A�je���L�d����V��2�?�s�0��)pA����i�a��2����w727��`�U�}�둩�*}�>��'ZXђ���.Jb+H�vr$���߭��:b71�4���;��:w�Ȓ���-KW��Ä�ᜃ�@�8���o��1y��`8�
��?RĆ�c���9o\��Ϭ��d�u6t�f�2��0R�,��f���9s{���n�
��F:*�����x�5e�-Z���W�	'��]R�������x`*�քS9���
�G0�u�\�Z��MdZO��ǿJ^��WAUK�ݖPR����tD�0@�џ[0�j��a��y-�-	-�
�A��Ŀ���a�p5.�d=���#�h���Jl�A�vf��H\�4��AI�������Q����n��0��~�b���`S�Iz����2�|���)G���j7�c��o�8$�Ş�/ޛ��Z68����5�������'m�t�s���Q�F�t�5�W�� 8G�/P��\��pOH׿����q?3m���ec�0H�+�(#�1�a�o~Y<�s��v?��Ý0�k�s\�<��_�P�D��I���~�5�mB�~��Z�K̅��(�����l�_�ǑQ�L4{!��&w��F,�[�4��)R��n�/2�c�5#�P�$����l�x�(��c96(��A�B)�^�;'LxI�M��݅�6�l��lY+l����\�(X��@lƓ��������k�'�O�aS�`@�-.heoJ������Ί�X��Uåo�����(2��ܘ`G�5ę��JrV,�O��s���Y��I�y��d����)��*���)@ P�@-����4�F�g3qXt�w���c�0%-�E��4�d/;�O�:K ��qK�~�-6D/l�u���xa��8�j�0���M�Hx�xq��T�a3��2!���.���ԥ��7ùz�ÄL��ȡ�����G��#W�Af�أz�n̦}3�S`[�]��O���C�ߢ��Qs�!�JT��ύ�=���������h�<��s��J�n� S|1�NP#�d�ǸTB"#^����N��&��~��#��v�5�CϛbQ-.�\ßM�}�(��M"oȮ�,A�*�����rbJ�V6���<�ҩ��;u��/�S_�Z/ཤ/�0+d�Q�t��,Yv* ̕=`���J�NU��y��kD�~H�{�>r[�%TV��p':�͒�;(Bj@���4u9��#@��o[$qP.��A�ܱ�$��{�s5���������#�a� u���	����f�cL�AW����<����`D���(���ؔ�x�4�Z�|�1�P����:>�,�5U"&�u�f����/���әNh���v`;��q�1e��E � e�vٿ��F	��8$.a\�� w�=�=)��?� ��������Nf������'Jj���˚�ਫ�@f��+�� �E��Nkm�߀QM��D�pM�M	�բ��en{����l�ݿ�����"�a�����ܗ$���_3bH�WfD�Os�4i"Ծ��`� ��Xd�U����x�}��+q7�Q�
ASY����s溶et�t;��S�x�cRU)�2;�o�q�E��۞�6.��ϝB�����4smM$��ӎ�^��m�W[�J%�b��q�w�=��q�V!�i8�J�<	�o+�0�T�g������ ��`���Ɔ�m�*�x�p�G
����$��u.��M Le��ӏ�����T���'RO��Pa;�ڬ=�K'�r}y/T��B��S�F��o��ժ$G�TN��9Q��z�D�xG�Wk��R-��jO�]����PG�.pE�'�np�kA*M4�h������3e	���}���`�"[] �S��;&
�iW��)��n����2Ԗ&�y-��ȸuS@���/�챓Gb<Q㷢t'j&��͍��-��z�	9:��6槭x�H!���U���{��:�-��)>q��=�*�c՟�3�^~�|��Q6%�"����4��N� C��9�ȫ�a�����Z�C�J0����rɪ��W����zڙ��5��f�G�����vnFl�1x%%�Ɔ�#�o���ח�3��H��_��T���Ģ�_�P8ŏ�z�A�`�a��Ԫ�&��j���X��YGI�r�(ו�q��鷫9-}�(=���[
e� b�ҩ4����h����(o�Ǎ��������oq���ԋ�����:����$qD���ޞ����_�l��S���.Z]2�����q�!A"%/�e�}�}rB_�ݻ;�m�?"9�Nɧ��4�����-cteP���9�_<=SEyV���Nل6�3�E��L%7`m��6yO�vK�f����k�txo�秼���2b�} +l�-�`�� �)^�@��I>͛�(�`�����؉�=?���f�����%P�'=ԫ8����I��]�QNA@�,�b��1�a��Ł�A@ɝ��!��Nv?�,�Ӯ�E)��ا�p=h��E�����xX���ᢂb��U�cDsyB�u�7�L@�L�ȯ����u�_[��4���u�q%��_6�g�Uk����U��f|�g���y�:(�6�j����}{�:[筍�<l�T�a���@���׽�ˇ�<AR�⒇��Y��Q(�jc�<ZO�����]'���h�\e�����Q�X��0{CAPQ$~�O�5�7c��b=�{
��k������Ⰷ�i�&8,�y0QIrA���}��v.�<C�.ߑ/��D�)�β#�n��M�d�)��on�֏��e��5��#����xN�ta�6�����W�n�M�8Cl����y$���RZ@��tu�"ROC�u�=��N(㏩s�����V{׶؞#0Jn�f���?�����)��ј�ޯ�	Sb�Ѯtk:
�'>��0KOnL��a�Z��2����ʶ��Dd�&xW�L]���t��\��uR�PM���혪�Fc�Sg�o--ڢ�0��v��dGoM��v��6�+�]	�^,H0��|R�YI��^�t���	��v5��{�W3�⽫�o*�g��Z�m'���Ba�t�9u���2n��;���7�3����υW�F�$fU�Z?�2��S/��?g�����	yq��mG�A�L7���AP)_��:>���j� "?��F�{'`��%M�/Y�[-�c��0�w�p)�Va2\Ք���?7�$f{��n���cP7M��N�R̤]�����r4�ڝ�_L�a_�p.��9hh����|~b�itZ��jx p1��������3<�5��#'��Ȭ�"�ȃ.�0[N��.�����'�ӹ7����@���R���:��w;��x�G��'=W�����d��kyk���p�M�2��>�, �bZE8y���[�1�<���)������S2o\N	w�It�e8,KG۱���'.��]�5�,��=�������X�K*���I��n2��Fڴn�� ��T��:�m�=ۙ��@����%V,��D4ѭ�gqnxB>,!�:�u9��N���q֗�k�$s��J����`]��I *g�/);����x�O\�R7e-_o�!N������x��q��G��u�t�&�B��}p8<��>�¡�ƈtG����j8�7�����(D��`0��2:$��WNϞ��}7O(���(1�"���Q��p�})������t� y��\Okk��]������w�o,���h��ׇ� �� feG���emV��m��۞�w������%�r������M��H9ɯ:��"y��[G�:�J�#m<��r��g9�����X
���!��^��֜��Xo�BV6�3���?��B�\�&�����P�5@�HOη�,D
���&�2�s_��"v0J(���Ǉ��B�v�@_jl!�r�\ңL�n`q28F�|�bK�b�t���q�3Ji.AX$$���+/�ox�FI��Q�.��5�i�1[!瘚3��/�~��1rL��-.��VSR�̃+�QvTǜ����wdg$h�+0�'�3{;cudG�e{G@Nm����A�=+��7��S�>����=5)/�����������09��՗
y#��QRE���Ν哟(���vXq�$t���$�Y�Z�go`$��L���_�:[��Ƹ�U��,�(
���W���j�%={�d��1���;��#��(�SO�N ��!��xh���L�����{�j/��E�#L&����x���Ve�<�8�ECd��#F��y�����I���x��U����!��.V&Qh6"�)���":��W�]xp��.��1���zU��r{1�7j}F궷�Z�m���N//̚P��h�����AKa�dV��&�מ3���R��lw��ލ�ë�؉Ȣ>F?����(�~ �`��Oٿ2��6�~:0�`�6�҃ق��s�r��~�HpqQ�������B�n-��G�������p�������0N2��� y��Q�ԇr�{5OLɄ��yȎO�q�n�L��:�@2]�گ6�u�B���j_ �j��u^ϋ�R��Z�BC�vz��[�~�;�S���29�T�6zS��mѮ�fT�X�.@p�b�c	�k���x0��=�Op �����y�������LY��cX{�[}@������6���|�S�]$㬧/:ʣ��Ъ�p��{�sBz�Zv��p�����O� �m.i/����r�D;�0��&�u�m�y(6˥z���)S>�HsAp\��,�9O�����m`�/��L/�v^� W�(i,*�$h���+���>W# O����I��_H���I���RIz%��Ɋ՗R�{��9�������8�!������v�u"�[��_�zA�xT"�r�ڹw�0).�J��C�3��8Y�7!�cF��0XM�K3�Jdk�t��$�x�;�PV��{U�G�B7�~Nnt�B ��F�>�71h>�M뀛���H���x�D��W��X�Ʉ���~��W�AK�tj�L��v��t�t��tm:�|�	��n����<���~�J����ɋ�<�>�z|Hi�+&�V"��S޷ba�hd���~&�s�v ȋ�G����^+ۉ	�����	](����"W
�c:��{JcG[c- ��  � �xF6
�d�����!�N~Y^��%�^A���*��P���#��ٗ�,�h�j�E��Q�4D��U�Kz��\P�J��5!�o�1d�L��Ni���`<�u-�߉Q'q�[�΂�Ŀ�,�q�4�e<?�����҉3#�v�Z�ͥ�}�P��e�S��S���1V)%y�w�^�)��B�iQK��*����
�cN����'���L�wro`�-�F����?N^n���'D�S�ݡ�GF+0��Z��Tү����~6S� ��3�wp/�R
�������y\�'F�2��eָ��r�?Z��	�F÷��5���}������j���7rF�a�`�4���ج����S����j����72����}T,55�)�Wq��zDCyq"nmh�#r�$�4���0���	R�Ԩ��RI���Z���`�q&<�lEg_�{ħ�B5u�v�]k^��j�P��#�l�S%�:���M���-���!�,V�$<��q4�R]zH{ė�B�]� �Cw����V�?�� x�wxd!�u{�q�h5��s��$��J&��zd�������`�l�!�WR��rX,�����$TM��U��̮���������m��1ɹ�r	�,	�x���`�ca���Yj��{T@�ϥ��t}�}�h�abڤ�s\h�TX11riI6R0'Vui�M�����&QvY��uT�*zw����{�������~٢��$�c���#�+�٣4l��tn�}ʃ���:���6v>xp�`R�QM�h��2��Q���l�>^�ˀ �o.��c����p�+7�(�{K�R�B�X�������Z����j�i�u�ם�#�Dʚ)8:&�=__�H6q�2�,8�[z�kƹ�/)ӈr�H��1ȤA�����������J����kZ������"��#�z���ʪ3��<q8L�zF�Y����D�����8}3ڈ�P;{��7ǵ��!"�n�F`�{(���P��o�����QԈ�*~43F�R*/B����~OA��}D{���	C����k��(��P咪��KNnyuV��/ �>������FI�O��V�8~���P�6j^���/�2&����&9�z�  n��h�Pԁ
w�F�K1�߸�P8�I�p;��ѩ�IZ�5�݉��~������2P|�~:����o��o/�o7
T���z��-U��rs�b�ˑ�p��a�����g�En�N�Q����͉�bF	���ĤMbD'f�@m�/Y���ѝ�bԘr��+��E��T֚P��'1�"�":����NKzf4:�fw��I��`����X�0q����ᖸ��'���P/fB�I5�����r�ŢJ��:2�|�������s3������ª:|����@6zR�L`|�Q�ϠѪ
���u�{}-ؓ5a-���y�ޫ�2w3��7Ӱ{�㓵�s�W�Gɮ�����Q_�R�o��r�h����5�~��K� EI^�4�Q�0\6��w(,t��0�$�C��_ƨ��ȱ�|����f�5x
ME��ն?h��k�!�fp	�
�H)�N�W�L���c(��6�-��'&�ҝX���@�_t��e�j�l�ɵ�E �����W���R��=�F�5�p�����(���Ѹ
J1�ڗ~�D�t䛡R�=��fC�4�l]����-���L�'s,^ڲk��� ���,$��@�� +Ru��� 8���0����s��>&��q$R�l.3[b�0	�h���:[̂kї���{�I�+��,��h�Hi^�0�^w���i��m���u�> W�����fd�!�Tr�*�!0�]h�b&	 �Z.��f���[�ؒ�|����^�v��O�@���EK?� H3���hƢB�����1�E�6�so|ꇧ�b;5�a+$��t5���{a�7rfJ~�Ev�Ϻ�ww�8=�@���������rBd�p����,Ԃ~1�0�UE����{d��V/��lbY�b7�iϡ�^�c䙌�U�^g��x��Q�o����K!,&@N��� ��_33m�u:�A'\�w͵ʏT�����n�yv�Ŋ�����I�EbǠ�ccS�� qV&NXq��<@�a?�l��>�}� V������m�b����X{��꠆��4��.6Z�N=Vܒ�[�[�@�6�FM��yo��_[Y-�ad�^*�~>��pc��3UG�֭[�uG�n�aXM�M=�mX�<���^��h�OJ����.�F�S�0��R��K��:z�)��ѽ�2��Nk��V��ʣnN�	�2�門�(MǙ�,��cqi��ىm!���F;'<s1�㏺sc��"-�b���{S���������:�E�v������ɠK�l��šc��ƻ��:�o^������ao�2N|��NlF�9�9��xb�y$%��r�e7���`�@1���RVeQ!�`�����فa�L�uE��HQڿ�Ѵ�|���V
e������u��K�m��c���G{Nt����A��tS��ی��/z������)�ئǑ��h���儃�Ƞx�,$ʊ������DŦ���{���	��ef�n%Z?��tF��B�b}�^!��!50k�曖��ſ-�}�`�k�U�:����\9F|�HN*����Ձ0��I	�?m��w�ƭ+�pO�0{*lu�P�����K���k��0��k��S��Cr6�)\"j�ň<B�%
5�����;��=���(�u՗ϞV������7\�؝�����鿍G�k�	cN-���FƤ�c�S���9.G@
j4�vEpF�HrQ93�GKZ��S�ݔW,��#�0������~ �oʼY�.'����� ���&�UX1W���q������(���Y���^���B����h]�<�#CT�_Y�K��TG骚�GH��J�N�D3�X������h��FZ����Q^"�t��Ӟ�Up�XH�ʸ?��Q�ţ&���6F���5Zǘ��r�x�M;���r��$�t0u��"�5F,��ɖDV�C䢡���_�w[C�u��ġ0��A�՜·��r�Z���v��o,@d ����s;�JJk��C�{�֛Â�#Y��9�E�o�YЩAT���~ȼ�{{��p���M�r?�Ɗ�����J #�PN�d�	RQ��G��3��}��B���������ƭ<["�%��	x;^E�ʉf�n�&�z,"�[)�9!�C�;���v�;��B]h�2�J�|Wq*���=A�
��T +撡�9y(_?��/M����R���;�8%�%dZ�~���Rh V����pvU����VW�U58�c�F�v�.M�^��ȉ}���u3��Q��٩��P\�%���p_�D PMA�y�n��w���+F��^���:`��I-7��V@������h�t��#A��$�y���L�
�33qQ���^�ߎ� Ze�9��1�fR�"��eۡ��49��
5�5-l�R�z�:g��iC�g�,�a;������Y�r��G��?o�<�Ttp=����A��y{`��J!�Ǹ`'aAX6�wD#��ދ�Az�IA�>)� ��P�%��� Bk��|ݖ:X����Y�)7�M�篏Kfe��� �k`w�=_����O�y��ᦔ����Ɵ i�+���E9�b�|�&�v²/l9�6���h��&S��,S�*׍�%	u�G�w��|�M�_!n��~D��Z�����Y�G�X�iC#�K�Ni�Yȫ�}�1ڿI��s��c��v
�l�L�6��V�C3����z%�?P������[���F��,&ո�SM���c[��\���PA[�&ƈo��WD�@��=��/��<��[�[ݏ��2�G���ɋTi�N3Nb�.|\�����\6��ވU(����Pk�+v��N%U�M����ؐs�H�/z��b�ךe��d� �a~á�?Ă�0Dde*�Z%���x� �_�m�q���¹����e�CMN|4������+]�z.���Q3���g:xΦ� �#�w
@}�P+BG�^�E$K�:��lݰ���$����CEw��t<9uTȷ��?��l\����$7��z���$<�d�6�ۨ����N˥dpNy��(D�ˁF�$:�����[xיm��B���ي�?��,�X�s�I�\�;�l����WK�Ċ��g]ɯp��ʥ8��0�a�u�x8�wgdFW�K�؈p��%>Ǝ0��FTq�R�~��'];c*���1�u��	�1c���p���k�<ni˵7�8��_��)�b�4/��!e��P�|A���;��l���8�F���ﳓ�� �c$���ZW��G��X��v�?G��r� �mg�)M�U�Y�Q��]�$8��ݬ�f�{4t¤�:<�/��|�r���g�_��₃����58���8||��w��'h�K��uҍ�9tЊ�,Oe��;�t���VA9�0􆯞_k+�����޼G�?d����P8@�N�'0ӁwO�?JƁEs�n*љ�[�p��Y�?�̃���-�g��7��#�=���ou(&��c��;�M��A��:wҽg�G�V�����7��3u
�q�ha鯜��J��x� G���ֆmL%�������4�4'e
Hk&��nҝ��
�j������t��7)&�;la�7�7eb՜R8����TF��X�O�ȩ��#�ni� �#6}�=@\
&�T�[��R���%3������>��-�=���I��/��(�8�2B'���є�-O˅�V����Xc���(��Qjx�XK^t��CR(�~�lU@Y�����n��o�g��{,9��O�@Tp�������$}|ϡ�%v/Ek�b��!^�@��� ,	Cs��W���!Ϛ�w������s~��;�і��+P���F��]�~�pV+�%� U��0DB!�t�~]��1+��w�u�mB�Z��􄣍��>�T��*�e1l����>Z�sB��wЋ3��z�ټ�U(��[�X�'sI�����~bx�*��Z�ȣm�f��j��i�W���5.�U;G�������]Ҁ��1xS���]���tmVoU@�:P@��ӟ�Дa�j.���\�x��u=����5-�	;+�ʉ-hRƀ���CZL{�p9���[��UA��7���J'9&��,��,��3��Q|ɤ��k�Ё��V�S��z��M�VEo:5�~Ӂ7����o�$��
|b�r�EƆ��r
!{�@bj���8m�c���`إ��zrK��|��_/��$�M����1sȌ�k��⌇��b��PGL������$����v�*�F�`jpn�S#��E\	8e��3�Jb�%�����q�~�?�XƟGL�7*�6�G�O�:9ɼ�����F���$�����qr[y��m��+J�\���[ں�,���HȞd)+�-v�s�;\�8m��m��1�9�.H'�ů3�^y^��$_'��~�Շ��d���:y�������tbƓ��؛��~��5]�M���?q��F2��y	gU�'�Fp:�O�w��QĴo��C�O)��[Q�pMS����f�1��)��I�����F0����m�YE�hcQ3��� h�c!�1����^0{S"A (�W����Ss��׵�u�	��Bs���5[�`�
�V�w}c~OE���G:/\QD�-}$��Z��M�?��y�G0�t�-#N���9ތar��xv�j5�����x��0@��"�m���S�1����0�� %�M&������X�Ry��J��^f�Ů�����c�KC�����^�t�&�<H�^R]���O.��e�j���NQ8�����B���r��
"�𥔇�����l�(	��������]����m��!#��5����u�����Yk��������싳�,�~:8�A��<����,�FN��k����O�jh1-��<x�+FK@5��^\�Tݕ���e��'�#8�ӡ�� �\-���	���@h�u�u����*��98O�j��4K��'�#��%S>�6q���ǥ�r���8~݄BՎO^G,s��O��Y��V1F8ٯ0�k$��H�S^۪���(U]d�m���-�%���A��eJS@�A������_J�1���P\��Ԟ5.�~u���/����)_��P��m�/�G����a!<���^��л�DD�߃��**f�����3z�5�h����0zw�/&,�x��B#��5��hf0��CUL���1���m��arx�r��d�F�  ���z��c��n��ɛ,�c���u���I�]�,��7Y:R�3%7�	TF���Izx���W7
W)m��3�]E������"�g���z�\���9G�E��?ESۓ�x��R��Z�đz��� ��F���~7�k��k�V���lr�oN�}[��4Ritx����t��k�z�+�ԩ5�#��0_܁e�S�/ɱ�D����E�P�re+�7�u8#�%G��#nRx�~�:ۛ���M��1�d��M�gY��XtU|x���*���%�U�,�j��ֱ���j�놅��E���\�o�//���4���e�����q���y+�L�iW-�?�|�0wrK�	��xI��z+Bo�Su*���A��-�XUA
co��
����R0�.[y��,�q���1��w^���qR��m&�@�Nf�E=,����U��aB�|+ZNd��f)�۱���ۇB"�ʵ	�
�N?k�=����${8��.x�t���#飡yؖL��~*�B]C��ׁ�n�)����{��&{I} �Ϡ�Y��2q�Û�L��_�DV�(*T�4��(I0�Q�AP�{)�s��<�X������C�i�)W!�����s�ʵ�ʂ��O�����2�e�2�м�ɟ�eF��{a�-�L���P+���ji1�͈������3@���S�TK�(pM��N
˂f .+?�4��_Զ2���J�.�y��G9q,�%�a)�k�<"q�nQD�V�dj��h�&�3P���q����_W�e��CRw+E�R|��Nf�o�cx��s6>��ib�G�-/��/B���gĘ�`���6���Z��@���jN���/Ё�Q)���
��p�E-	E��T�l����qί��ys��sh}�9�,��L��%�=��	�h0"B�0¼�{� C��8ԑ"�Jh�F��Ͱԡs����b�1���[$����� u
c�&jد��b�^)����Ș{�<|
���j(b{�� ��8�1[��_�@o�_'�-�����]Ӑ���vIV<7�R��^j��	@�
;�����R��ͅ��9��ו�;�)v�n+�7�ag�l3Afb���#h�]�1� ������K�%�\Ҡ�����3yO��yK,����ݱ��+����0ӥ$`�Y�/S��80�;x�(|�u�D�u�`�U{�J�w=A�I�&��W���Q�8�Gql�l�0�P��<� ���գH�K Vp/��ę���y�M��.�N��s�А������e��/6+�A�E��ϰyK���K��U�j�f>P�n�f�������N���`�MI�$i�mZ"w\4^R�ghlR��w(�($C�Z�ˇJ���=����ފ~`�s�W�zqH���'r������p@���?��pΛ���;$Ɇ�&~�T�NÛ�椃ߴ���@Au��>5��.o/�Շ������D1�ֳx��aѳ��m���r��/ɝ\`���%rzlͭ9?y���)ɭ�w��+,�:���Q����;L&�����\�i3'!�.�8WXs��b���P�{P�V�E�<yG�$ڷ�}�s��A�rS���u����Z����U�Aj�i�/1m�в�0qj�ϵ�auL��G�� ��`l��̶J�r=�,���^�I��o����:��J��s��t��C��p�(+^1�/]�,��ӄ&�|JOB���ﵣ4�(� ��I�p��,p؞����(��@�g&`"ԛ��H�݊�
l�(x���]8�������hC�C��y`������V%+�&��X�!{Vzj�Y�|���p���xb��:���v�,s�c���\{rU8*l�1���ĝ�mn͍��
��d�a&�9r���ئl%H���6/����M�U"
��H�I�$�e�h���嘲��t횵eF�F��V
�,D^��g�	�Ya�/���I�
gaU���Zt���މJ�)�����)�Ao��f�J	z���u�G�9|�I���ȸ˘o���*�x��gv�Ia��bT���J�g�my���n�������� ��
O!�|����߃%R$ӂaP�����=����6�T���A�)ʞ�F��Q�\�����"^(j"٩��2ڷ
<����h�],�u�$�_�5�{�d�m�Ȯ�ƚ}�I��bA���&2���c����'l�#z崀��Z�){pL��>x�Θ'�.fNd$��Xa�G%k����Kh���Yi»����r���>T3dݥG�����Y�G@����sP�ںÂ9�2�k5Ջؚ�>)G�j#}�zN���uH<L'���$8^n�{+�E�R��6p98V���kJ,0��Zv9�`y<����BN��A9t�v�n���oX��,L+�2�t�T h���X�Q'-H�%��X9'��0�G�
:����P�Mg�EZ�w��g�**�_@KG˓+�)8p�/��>�8���ÂD����yc
�$��g�j�_�����z]�i����@�ק���bH��=����u�'t��.=($YB�e���L�XY��X�P�&x����ܯ���,��#�2�?�-�I/.�8s�2���r����7���\0�W�gR�n7h
��˞�Ǫ!�LA���w��`�KFX���4���D*�i�X��-�x��3WH��������jSǷG��v�����탳�q��V�� #�kI���&h14���`j�j�·���U�.�m(@�N�EQ+J(<6ҕ
�;�M���Mo�� D!�x�j��1�]�Z�'߯�N{����F����5�INX`��7�݂��}���#7����)���:�(��� b%A<�u4�����BK�� ��f��c$d�#�&���n4��&�D�G�O�A�GfUr��9�r��h����� 	A��F����d��V�1�>9y^�L$�S	`�I�P;�0N����u��Q�z9��o8�e��˝��J��	Jt&������rܙ`����2��Q�!i�L��xC:�E�	�\�ڝJ�qV�&�]�x�J��f1Nw;����Y$�v3�"�,��MS�G(1�d�`}p F�Ǥ0M�L��A�&W��ﻢ�k6u�,ҋ��i�ɍ�>Ӗ#�X(]������(�7��@fG��U�ֺ��wR�p�X�s�j4,���Q��Jh� ��t���+$�I�ڂFʹ�v�X�T�3)B��h#�,����vo��ί`�+�o��n���]�;�+ve�<n��o��eX��n���.[��3%�2�0B�zD����{�z \��'�l?�uӰ%M�ٕ�h�vǲ`Kg?��
\T:�O�)�Վ)~��gyU���7o�>m��IQ��n�;���An�9���XIw���7y`Ne11�W��NW)?�3���	uP�$S�
�ޭ*����ͼ'�p�X4��jF������?���s�/u�{Yj��
Ӎ�}�J��̻�"�R�n(����٦<���x� ���g�Lأ1J��	�I�˚��e��(�����UY7�1�r+q�a�;��m����$�10�;�T�C,Aۊ�(�T��Z�Ҵ�3�'@��t/��w�GR��k��J��%�^l�|L��Aw �c_�бs%n�Jh��A=h�~yB������Dh?�|��h<��3%*���dR��m22v
֙~�F�<� ,�Xu���1�UIF��OT��%���P��'�Ճ�&_���*P:�Z뷴b�l=mH�:z�;@y_p6���Y�� *����p˒��)W�����A�d���� ����;�u#�{N�X��f�>ƞvpH�*�G:�#��)]ڱ������r��]$X�yAl�¢�A��65�K�0�S�K���[�~�J�Ќ�3�؋h�	������]z�(�p/"unT<�w�%a��W�L��FҨ����������>�L���~����F֍��]8�Z��yBdƀ��\��Pb4�a�E�x�b������2B���B��'2>�~2�t�"�_D�7�>��%����y�N��,�K�<�X����
W�?mk���"Ff䆧25��D��˳�6���A C�\+�@��q{!� �Չ�54s�"��0a��8�Q�y��k�����;AR�x��Q~�dx�e�mQ��l@�xL<F�0V��M�9��ͦ�V�:c	XK���%��?��|��&KLA��Ӿ�B��TՖ���� �Ӎ�A��I,�Yb�Ԣ�b�,��-{�LI�l��>�3}<�B�%:����+ȀPʜ�"
E�������ZD*K��$��ً�w]G�ކ�O�i(Hp�h�8�+�3@E6�l�X��0��  C_T�u(��`�#��a��Q�H�]8¨i�.!�=�lg�:;�&7�EˮGJ��2��:5��%c�Ҩ5�*�! bz�
�4ug&��8po�N�~P�?�_�s@9�y3.D�HH�gU9�
��t�;���(V��%%���J=��]�K5�r)G��\��[ƙ@�����{�C�Mpz�Zz5%�Dji_B��h�D>>�oEZ�/��C�D�edU����>��7DG��L��y�TO�{������+y��t%��c-;�6�c�#\��^�bM3{��-V5�S ��O�d�Z.�a��qM��&'�c�_y5E���e�� ����x��&��;���!�#��#c�~s5Tc⹶6��5�q�H�����GѴ��u��OY�����o���3��;TJ�ÛZ˰�l��̚� ��z��+�	��b2�s!vf�X��x��Yf�jSM���Q�ScIhS���r@�;$L���ʘߩ�؉���RpηI�4c��T$��Z$�rÅ����bK2�1<�g���l�x[�����ndB��dF�5���L��Ғ&�JwQr�:���D_�ɬ���*V����ܔ�2��"p�:�T좪�sz��B��~-�s�@��'d�3!����J�Z���O��V�(�f�4�ƨ��c�g�UN$�������,ckAV��>�;c�X�bn&�5eF�C�(�n�mM�\A9�]w���a�gOp�m�NN������ �
Rz��Rש�}<��[i��U��2q١Y�y��cW�#����6�(��9vJ���e����n��P�V��{�)����;٢�̮w�|�لԌ^���]��b�	z�1Mtm�s>jk�X{���T4��qF��4q�n4/�Q�CE����]	҄�ĉ�N	�T���t�w�u���m,��^
���t��� |����+ܲ%D��m�vX�:ٺ0�~�=�sI��jg׉O�9Q�'F]�G��9gW��cv����'�w<�V`��0QD�̲�Q���7my۹��[~��8(m��Ʊh���S��BmY+/��_7��p�,^����[��o,B.����8�sn��1e�Ѣt�u	�Z���w��dR~��^4T[�����h��)��� @�o��4����@��W��_�]���~*��׎GB��QQ/�#�3�v2v��6ȝ#�����Ⱎ�b>�Z!�_�/Fv�Y��ܧw}��y�$�����P>�����p�%���VE[��:��GS+�n5�$:�v�I�w�I�ԌN��g]��\���n�Xs�&���2����ަ�_�ٺ�Z�3����z����GȔ��.�f%O=�l���ZQd	#��{�% �P��5x�����vo��z��c/�*��W�r�/
����l���m`�Q��V�gl�i�.t!��%~���`D�H�ӯi�u*+]�T"�G鈣`���C+�[gg�����t����_��k�~���8&��b�*�����6�����L��L���8�7&�|)�4��Jk��1��%FՀTF��[o�P�V��k��j��7��V�O41�Flކi��(�ץ-#o��Ѱd������W������ؖ�H�{�iP!R�.����ʮ�JҿY��2�T������.��`��y���� ��=�c cQ�o��S�%0�d�V�ܿ�	��@A@����DU�LUn�A1�;ۉH�@����oA��ޓ�k5F��ق:�l*kj���MK�Q�+��+X �x���B�\��p��԰�uA������c%��{��Y�"\�}�n�9B)+�d���%�d1�ꐢ/���n��\Ю$�Q"5�A�fĐ�_��ο��ڟw7���g�fX�\���C��]� ��w>��_:�t���QȮ��.�|�@��J!l?��
�"����]�_Bϑ��rk�\>}�7���,(W�BzZ��g�6?1t-�[��d@s´��}Y��q�_J���%����ӓ���搅��k@�"���2��ؕ��s�39���5X,�hj���.�b�����K-K�^�l'�	@�a�=���Yӳ�>CXv�@۝LHj2F$�y`�g����nEZDg��*���~�y�a0��#
�&x����x�Z��[��9�e+M|�k)���-ٱ3�vD�M�O�0���5�7��~�����r�#qf��Z��֔�H(wË*�k*%��:FɰJR�D�MA	\� �|:������e�G��eЃ&�?���m��'�8+��Y�w��m��L޹=�m�\�¥QP�v�)����;��>��^[/�&ףZ�{(5��-W�>N����"�P=[f����=�o:
K��ٗCE�y;ax; G�@ ��a�S]݅E��R
�^B�Z���0���Z�R�F���jĴTir�F�����>��Gb�2�?$+͌
�l�Ӿ��!>�6Q�V�1�L#n�6�؈#a7��cz��zBo5�>������BpC�@�*�M�1���,t9Jtb���ɝ#�G!Gz?l�X]dF� �n{�.pz}}0���s�������G0��<��6�j�[��*� �A��'�b$��B���HKK֠+�z���!`+z���$�_�R'F�oX4`�f
��Bw<����q����P$����޿���$�"�L�u���QX� q��<�*R�p���K������LOӕ�4uP �&.1F���H+��`�OLl�Su'O���c����"�F�Mג.� ��E:�'�d� ���VK�O�ױS��j���l��l�v'�� 3���D5��臨��@N�C�7�#a�sh)S\5]��GicTmY9�.$ńM*~�-$�U}�!�G�z@�l� ���z�ݬBed�����\�EE��Z�r�ذ����N�yL*�;�@�GP�E�vA�8'����ЍD�[�1S��9�5i���+�"_6j���$�A�mB��Z`	���Ve!1���wV2 zW��lT�����*߅﫩��_��i��l�,O���}����s�cN_1U^����`N=#"�P��K����.����q�~���nuy��'��&�u���	�wF�m�uo\f����+G&�_m?(����]���a1�=�D�ܶ���ϒ^��xo=��^��iD��.��v�=}
����y ���گ|�
�$d[	���s&���˛���۪󪺽�~��x��������~�o�����z�hnQ9�jn;e�0D����>��d8��P9X�j�����Se����ZCJ��j�<�v&���T٘���C6Y2}����"M�1�g��8}�I�g�X�n像��) ��	�hG��_Ϟ��6�d��I�.O}`W��Ks�y�9l������k�~�k�5���o��}(8ݩ"��wr������ڊ%�E���Z?rZ����j��V��Q7���C�z�����|\�_N�v,
��vS�j��ɅA�(B?�����aIA�oT�Ko�}x����\7�L�aY��
C&F�Qb)d��� ��c�L��=�zaN�x�5P�=_K?�G<ZZ�YL	5��WZ�&D��4�
�D�U��ůX4-A/��Ow�'��l
����<΅N����P�c}���R�ԕK"��"S�>VXB�o�ˡW���$��_T�CʪI"�ǌ�n��ݳ���VV�n�>�+�?֜�sl!�����s jW/�w�*y7M}���3��/'_`���8��!(P`�A�T�(�]����X����8�+���N+���p	V��ԕ��5\9�)_�ھ2�Z�'��J�r$�d�Q4��.�%AP��삟�PP���R���"��2}]������&���N�m�.TQ�B�I�4�ȗ�a��7=����M��{s"���E�)���&�P�B9��Mf-X�蚎����`=h�6��|R�#���]�><	�D����r�������$��1�zZ��-������^���B�՗���*���`�U�壕�V���{�@�^�Z���EI�8�Y�s�O_��}ǭ�3�Uއ,��B�p'2qZ{�(kb����|ئ'���u����_&���*��=3�ѧ�W.>
�4k|��Z�1q�7y
��U>��+2�7(��v��d{}�(�&��XTU�����D����.�����P����Cy�X���&�%�W
�:\7 ��T"S�q�0R�?,f&)9#�A�O9��Dƌ���M�ްNϪWQ���-�������2?�L�a[K���G�SPP=�;�i� �ʚ���XF;�a���2��0yYFS�^�!��{�7����2m����.���f������bX�Z>Ŵ3S�mFS퍟W��VW���WI�e����AFm �Fo�e��.�X�jf������4,C5ԭ?�L�������9��x�wE�A�A��Kl/�7��-PO��F<~��G���M��H��JF`�i�[0ıAq�H�@3������=A��hE��ŷ��#��k��X�p�b>��D�F��l'�}��,�,pv);�r�w�u^���l8�y�h=�`����޳��.m��%ȰQ�&�[`$L�UM}o)/wW~!� �QB��Jm��	��t��s(��4�Q᠙�V��*[��z�ƽ���f1ǫ��Rh]?�),!򨠊c�GBT��+���q/�Ⱥё��G͕ƙa%�%�#{� &,2)�z�@q���S�8@�wN8��y����^�أ��ÐoI�:�d���j��-�q#�a��k���:�,�W@Py����{ F�	�����%�����0v���s�����a��
:���-}DDl��?�~���r�Ѫ0tˋR��򿰲)�|�loGP�w"3M	�O8ˬX{>��ߥ��7O^w�KL�E�����w��|�M���ޡ2o��^q��H��9@�ǵo1�9�>	sY:L|_4]$Γ	�s��� �9W���O_�C���0�����RI�U�m�7�;�+��g�e��o��ê&'������Y��H�؀�4�ʘ���Jތ�a�P<>��b����ˎ��J�Ι�v�?��e3أ���=���aM����[���F��O�K`(�tm7�\q��h�/(�H�y�#��k�f���;v��%����g��~F�!a
�l�$!�b���^t�o?o�3��'1J)y�l��قg�-����y{��<�+]d���a@_���I���[��3Ny��T������,���%���N�Ot��9d�qͽYS����M����{&�})�`��:O�g�a�KuQ�2Q��o�<�կ�M�����3^��3�	z:�}�/9���pm^�v\X�������KB`�K���1�M8��oj֏_�����
*z��g�����H�?����yIM��Z�	:'bX��IB�,�?��[=�"�Z�7���_$�FB�yl*�~�F���~�A �����"1kږN�����F���|����x�Ud�x��J�D�}ҙ�<���� 8r��1�����p�I*x
C$�!+�K�'R�taT��K���)I��-���N��I����A,��AP�|S��9^��R���o�}�$�+m���|�n�:nd�A�=�D�Q��Ȼ�!a��(*��zG	�pyX�Ҡ�I���gm�x%�8~�>
��1��	�d�ПR&���+��4�N�-�T}����:O�zG�f�[)�F�
����(�z4��I)�N>gi��TgFq���N
qS-�R��C�Pi��~Iw}�*�D��;�����yQ�y�'�Y�	�r���1�{��S��O"s�9z�l�HIM��1Â�6bd��S�j�нs)�+�'�N���h��rl����<�L��I�.\I*���fI����Ng���BO���KNh�D�ZÊ%�߽�-�F`��v��S1�dT��I� �}���)�`g��x�a�\$cu�vʵ�Ý��O����HJ��[�h�h�
�0�/�o��K�t｝���{M�=��3C�7�.�cT��9�v�,��t|�)5���}�?��3�K>���k(��ol�{��l`�lL�z����7Ç�߫�^����Ͱ#�Uh&��[�ߋM���4�;��$�lM�hF�qF�Le��d�Y��خ��U\*����& �J!ׄE�@�c^�qSՉH���aՀ�Fݦ�VCd"N	�f��j��6�,D9fƀt�U����������7$/�gP��$%��T�<�6ؠ�c��N�Xa$�r��˼%
{~�y�)C�!Iw��k:�L���*B�T�U�1��?SК�]�t<�> �k�T�]�CT\Pi ��6�)Th��S�зmWp��*���-Zε��L`lU�pT-;��'Gs���6VnD�*wV"8�	�aS��L:��RVeS0 π��x�o��=i�����S�ܚ�@����p��Q3C�f���,��咽��7�y�d�Õ��:�^^��X�C�L�6M��Fo��jeSY�W�ƅ�M2&��9��� ѕ��zt�]���������tM
8��T@�V�DGy�*�t�w|�dg���S%G4O��R����1��2Bՠ*�Eן�^ξ�����{�����R�dn��l�U��GxW�L�W�%W�,����d؞�J��%k��-�E񐛿M�a�U�Qx�PX;CQ��Wb�"0� ms�g���Z�[�~�R4���)��0q)<����1� ��"����&U��K�|'�`�Ha���7#��g����v���*p?����\��=k����O[p�Rwr"���*$ JU�v���J��0���EoE�%�x�������e��Ф���ڑ�g�6�+��Hr��h��\���+1�`��K������"S=��ļ���j��9 ѴXzb��N����eMsq��'��`��8��+�JR��D��\�� W��Y��!�5浟��:�*�{L`�߆pG]v k:7+�±�����ǖYƸ������	mIn��^ŵ�|[�[����Δc�,¾��������~��kxf �G�0�a�s"���������U���U�.��5�����}�th@Q�����@�8��F_?~��CZ%Ưq�ѩ^�vɐ����9JԵ��ӵk8�E�jG�t:c �԰�T�{��}<�s�QՎ�ٚX�d�
����V`����� =��S�Wx�d�r��S��������i YXCϰ��9N����&�N$47j�(��!�\M>}���q#���,�&����0Ŝ��h�.�z]8�NƟ��{.�CN��'&��*�\p���B@�����߭���rt��!� #�6ola�C���:�|wE=��O��-��z㽁��W�����N�`�U3���|,���a|Py\)���HH������ETCa"ehr���buٜ O&NM�||9��m������G�r��_@�j�'󀼐��-�J��O��n�Ճ(�e�|�au��:#i�{�bE��:�b6!ME/��q�J�*�k;P��=~h�'��AF����͚#�w���z��
 I�m��9:�(b�P�{��k��Z�d�*�RT�W�P�	�&q�A�3�߬�7U8�GM��zslײ������34�>�̽e��"�����!+���1L��'��ٟ6�a��*�wR� ��4
��m_�`�������~W�zQN��#��"����	?^s���Hn=4�!�s��*3�r�Z���$L�V���r˘M9	�C��^��-����D��;�eo 9e$:�{��m ���k����~�>($.��9�	�K�ek��?�,ٜn�a_F8��	�!���Z�bS9-b92��VTV�*
�j=�H�V@��J��> _�0x�q��Q�D���X�s�-��p��X8�Ѫ��\�	�14�O�2FDZo��-�|/�
�N��ac�q����^/�.�;�|VL��q����wo?��:�v�CO>2.�H���q�n�-gB�������){����EJ���d� �B�@G��K�����wdY]B��[Aė,a6/�*��|D�M)�ȯ�d�h��	�!!>��z��uC����؝dT�a���R�]q����8L�F�(�!ȹ���<��Й���c����eY�'v����Ijhv9+J�0��l�*/s����J~�m�@��s�FIe��*�T�ܤ���*���'ݲ\w"���P�s�i$�q�}�eU_���������99�<�*� 9P9�pEW�U]&|���S^���V���^���ݬ1��r��Ȫ��|.��������hD�:�ѡ�Z�,�����7��b�',������LUF�`&"۽R\��7�2(���ω�Nƽ"0���o��t�t�h��>IR�!�"�=�d�m�j�1)��t���7�ܾ
U�K��w�wT��t|�e���D>�_��+�_��ڝ)E�x��Hң�6�����ì��/�Ii��P�n��ny�h}-�p9�<�(�R�&��sp\�:6i�H����M=T�_�~�aD�L��7�&��M��MP�zz��y6Ry k��d$�.p�Ն�6� ڈ���F1���0+L GӤ�c����D�� 7�AI�����`ҳ��&0lX��.��2-V�SU{leS�?Е5|Vp�U D\? g�Ѹ�ɓ�� \e��r�=�)��
rh��Q��3*�Ce���M���r�(�z5v��;�
,-\$���H�/����[������/@����Xa�[���b%�]N�S��P�CN��[���F���f�O��4��k\-1u���Y�/a(K/��r���%�@������m͍�u�a��Fn*V������_��f��\}�U�9K��X�P�c�S[�1E��5�Pl��1��H�o���ܬG�ֆh��S}Χ%�rWc�]�N-tWA3}A��ng��Pn&������ې,8��I�S�_8J�S���E�ՐIGÈ�\a�@3����u�X���NPd�0~��E!�|�^3�u,��]��ԉ��ⰱ�KM�����:9�2�
H��_�&�\0�5O1���^�FCH�")��M�w�U�)v��>���E�����J	�bQ�^�ȰZi�҅mV��8�:f��o�켓�T�^�4wN�$#�g~�]��<�&��eDI���K��@�IA�9����͵d}�����z���E�8U!�����:i7���W�}M.p�+��|U*9Ǎ�Q�8�4C�r�ih� ���5r�T�[y]$���_bq1�52W�L����K����R8� ���/���6����	��̟�����/&�;�r�
]MfwL����͍�t�i�G����¥<r��P�R>.���!�F<.ogɗ�X��{>?���t^v�T����z��o�������m�P����U�VG�
�Xrd���Ҙf�/�������x��3�Sz-xm�#_AOA`���!S�vF��y~�[��f�	Wn!#�>Ư=2���� �uY򬫪Ñ����_��M�z�"b�Uc�-ނ������ɩ}��x!�'ϡ
�{B��n����ef�_͖�U�[��Mf=F��M5���\�H."8��Er��v��@�҄��WLkN1�)@2��E\K�,��N�o
�t���{HԎ�~W�D�M��ޤsK�qQoM��Oժ�컠��s�M����^T�j�!`^�ņD7�zĿ�K#���Oy��R��>�wp���r��5v��z[��2���媙���1C�7ԣ�e�_�o�v19C��S���zܯ]/��J3��� ��im�]�?�ɕ4ϖ~�M����[�K3T��K�DJ��x�T6��ϩPQ�+ڬ�&���%�����w�㒻��b*X�;:�}R�h����W�F|��I�jӕaE���8�AM�����oۻV��Oخ��RB���Ư������f���q0��A`4ȱ��I��)H?_'q��2�.��#� CXܒ5 �.w\)����Z<�HkZ���y�_{�go>r��"�B��=�g<}4f�8~��9���uqC�ΙB}MH �O��P]�2���c���3:=7+ɍ�ϕ��u�=,���@��_@�b��{e$�F��TB��@O�-�8�.ڔ�U���S��}�v>D{�g��6�"4�=�k�ɫ�({��zh(n�\]�(�%.S�pz�m��uD�aH�?��M�P��K)��˾����ʀ}h̎&����?!oU[&���4Ϸ7�@�%�l奉6b��5�׳^�X�]���X64̌��^	��]q�ʞA��=�w�(�ĢoT2�@��5L+k��o�V蠬G��T�E�����,�4��VEwPI�A�������O�F������m�� �GH�eo�/X�zv��t�K�y|{C�"xR�G�&L��?5+�8�{�V��Xw��8-A��Iq��>��d� "�exc'��WlX�xܰ�B]{@R����h��A����n�@��+�*h��IzL�"���QPc��ى����΀��n��ڊd/*-��eKǙdf��dq���>��l�Vݛ~)G�_?�v	���?5:����^�J�q�$��n�V��Z ���\�hQ�;����r[� �	>3;�5�1j����Ͻ�U<�;`q
M�t�s&9_n)���ve��)�|m]J?g�N��&�%���V3R���R*Afn:)J��q������c�9'4��	y�Z}\�p���/!�� �dX���S�I�)&�U�W�kS���Y�1>�Dg[=��Jk�]_�2xF��Z�-��1�ݳeO2M"L���B���9�c�N���!��(8��v����FYc��$k��}��e
t�o�&F�������!����~�̷�كgᒏ�_�?�-����!�s�!ytp�.��Rx���)Q.k�?8��ڀ�ىa�\�W�ʮ�{�Y0���@��"P��ږ�l]���]�k@�������J���
�]��QFǼ¸�
my�"�/
B�K� [����w�LGo������-��WSb��7[���f�D	|ey��y@�pN1~;b������n��0��l] ��AE�r���4��`�(����!�,�d����n�DgoJ��h[tn�	Cw��Ų�!'¶��a:fĳ�m�U��E�|Ly����s�-���AI
�ys#^�����?��?��mW��+24hM�1>W�q�lhH��@F��,���M{.����#2p}��u�t!H�7��4W��%�r��͹�8�|{����g�Ş�����UkH�Y��n	�7{�C�g�i閱T�l{N�=�X;}���u�ؽB��~̄#�xav�su��LQ'�E���I����tQ�v�C_�'�œ��%��[`0\+�C�o�D|\!"5-y�kjNe��`�v3^�G24�=#ͧ���E"���R��м�)�nh�7������ �_D��3b�0<��n��_����G嵹p?�� �C�{ ywE�k3(kR�GH��A^��A����ya�._Ba>Z�B��v�7X����-,�1��)O�)e50c���1QtK��q3�^�tyx�����jJ�@�;)xg������MI�G��=t�4]r	����(G�I9��f�/�ګ�z8x�G�"�kg�;���+]F�ǡz����_��>�yk���0�mxZ~�Zid�o%�?�փ^��4���D��Ea�1ҝ���v���Ջ&�E�q
Q�����F=5����\I�ɜ���g3범�W��#4��.�xO����b�_m�Y�c|{���&.���[�$d�!��1gc��E�R��]��)�(Z#��H\W��!7J�6z��4��
��\M*:�q*�KX組��Z��f��<�������$��Bh�,�B>!��1� ��NF�/`ɤ��C�%*�MS5����l~�7f���p%�T���^�{�����|O��%2߁ú�!�:Lv��mY�������;�D��p�
 ��Kw��Fһ��5��^�����
���q���Ĺ��7����c��ׄ_�7�4���[HI��x
�g�b�`��ׅK�3��"�Y���� PU�~^���b׺��8htx�y� n˃9�����c�)�0��[�@'#��MH�L�z��]��r_G�	"%�=D��s��{��$���M�)���\{�6ʠ�4�*�5Rٷr0�f��P��#�y�1U����j$C+a��T�e ��d4;�>�ɼ����V���BI��$^�Tє��r��p����!�m�<JK���m�8���{t���sJ�Rg>���^��+K^�#��p��[~��{��ͬ�n�݋��c��|��0T�����A����ӧ� ��߶���0|yOT�Rp�Y���������2��l�z�ź\�-���p�&�=Գ�#���%��G_�@n�]��@Ώ7�ۚ�K*�����r�m�ɀҷ
�d��B����j���e��)�"K���\V,�6�y��~L�����z&����~@�u���=�t�z9��<�b��0���&�����9㴀fRD��[?�>G��	�9�è&t�OF>L;���I���E~�p1�~�<���^u�V&8�%K�f�D���0��ZĦR�pB�ۈ���?��2��e�V%�CP���>L]I��$�v47w�7���BB�9��U�v�2T&�^˗r�L�c���%�@�B�6h��H�"�y�a"���Q5��-�	��B��!˕'é�L�hw�J�iׁ@�O��NݧA�,SW���H>�ٙ_��m�Ƶ���@~E��F�h����A�h�T�{+�T�z�=m�(�ڑ3#h����1m��V����$�_m���Mm\M����f��܇�j����\����"JA��g�ql��Xr#�醌E��֍fg=��ie8<5+�Yp(B�?�!�#��ps���j�8)���*Wyusן���c�+qs����lk�F�I��r���|?�.��� �͊e|O����0���[�/���P�b�} Z��.�};������D8~#�G���kgq�Q�I�a��NW�T
2
?i)��=�����I	ѩ���;�',*�br��z����A�ڻ<��{x�1��ɱ&�^1�[���X>�T��k��֜a�4�Z Y�8ޒ?�[u�rDaҲ��_OR�o흄5���a�,���G.)���U�'�7�K��)���������N���<z�4�i#�{�_�+��"aG����5*mJWjjW:�O�(�pe�:��66D^�o�9��dX}u�`��&/����[N����p��'Q 獐*�T�I�>=����ߐQL�B&�����"M|� }�.p[�ѻ��?2e�����N�Al��t��S��uwQ��D��e:�2��5��W|����}O��k���s�k����-�s�XMT@�Q�̺�����wzx�h-M�j�,wL����\A�\��nD��o\��;��(������� ��ψ[���I8$�7�&<︟�OO1؀��X����}�q��uM��.�����J�~��sX�����<1�vl��Q��$�,	2�=���m��o:��d�S �L~�����=��"W�.���ۅDk�F�*�+�06<b|h-��.C�^�I�*�4���IO>4���F=��Ç>y,/q̸iݲ�@��&�R�̤���� ?X�$������)E�x��E�B���mO�����zS�H����DS ee4�!��s-���p��x��F͵�h��M�[sx�5�!.�93��0NdPra�M�C5��XA=���_B2��W��)���&x�@��Y;�	��ٔ��}��F������a�h^�pA�����lƎ�#��L�+ �{
A����m�܏�Mj�/D@�6�M��D�Y������&9����*|-��'��yD>��y�/@���!8��T����mS؜�0�M�J�]<S,���w��5?��2ڠ�h&e����3No���Z�H�B:�����
u��,oD�%@Y{��A\�9`=N�~���(rB�Qn��uuBǐ�7���BbI:Uƾ����1kYg_���g2?c�k�9��f�I�Z��l��n��qqB��B�(��y����Uc=�6�!bn�5C�~Kl��E�눖��N�~���Ҧ�J�&�)��J�k{iSC���Lluڏ?,�:3���2VM�:wW�`*��I�_([�B{��A&�-5�vT�M�C<�u~4bXeCU��V��a�ແi8p/�����k�l�̿�\��Ԣ	�M�V�~�<c�h+��{����Q��za̗� ��۔�1[3��i��`2Ի>�#��>
~�iP�+p�)�r�]�T�g_���O�˷��/��@��Im�+4�a�Jz�蛘1kXG��w�Zr ���w���C���M����2�n�}�����@>�b�m����<>�B/5��#_�7�l�k��
e*ⵁ+������%FCq���8�22�
��	�c*��~�s{��.BG���<t�kdڢ�rda^��@�"~�Y=^�M��u�"�%�s;�u])g߼�nr�I{VLd0^�LQ����KH��#�*	�W�-��o5���c�&w�{�=̍֎��tX�4m��`�%���hh�>�/գ������d[���JF�JJү�z\9׮M��2�$��rz�9 `w�\��Nk��N�V��:"�ԛ����3sY=la�\a�U�L��D�� �%0j%;�%^�}/��l�8n����8�����~HE���@�[������'0�Dq9�!�)n덄�7n���U^Z�J.��-�f�y��'E�/�]���_j��G"ͫ�"t�Kμ��c]�V�5�m��>�ӠMm�z�}���x� ��iߋ��cX����_�g+����.�#��{�ה�Q���v�Oa� ��-�H��O��ns[��<&�����@�x��\�U7cx���\o�B��
�U��.��hL�C\���u6�ŵ@ݠ��\&��T�쩠�u ���u5m��h/iEąi����R? `�J��9�e<s8�s�Pt�|,^�p�R�g��\/�]vs���4C飝�k�E�%b�B� �N��Y�: F�AWdi�6��{�V9Osv��_z�%`�@���-$*6���)Q��2��/
X�T�<���b�3\�n����of�
	=���9��"V"-���/\/;��&�4��Ŵ���?Z��,dA�x��Y�8�l��F���g^��Jk�{�[�F��k�[���A�,�A�:��|���B6t�3C�W�s6�iB���Ow ��kB��Q?�|t1���z;Xz�i�L�/��@�L�c:3����2v��^ @�D�����N�1`\��`������j5^A�0ccn|B�	^t����X�e�[�8]�<��8p�X3�D�bp�b�ڧ��܀<E���'��q�b�6��XQ"Ad�g4��W��֑�~�D�<;^�t����X�g��R�؆qF!��C���+�]�`��.'{_U	{�Kr[jM���Jc�?�d�8��)�U(zKVt�J[+2|�W�N ��mj�$�X"��cO��z��+��q���ʕ����7)�0�檴L�j}�&!o{�����ۼ��t/�a��|L�'���Yj��(��A��%g��ʲ��_�����G�@_�"�,w8��W{L�q	����V<j齱��ݛ��#���#N��۳E@���w���0��Nv�Z��U|}�ھ���TnX�35�{w��s>��B�J�O'�"M�����Mn�d W�'Sw�&�4)�`��t8S�gr�T8�E�����jd�8�冲���̨�<�&]%�)�fj'xӈa�ic�����Z����%�_�*�C���DHQ��:n�f*q-���^�7W1�6n)w�J6�X|,(X�gÇ&���q�@l�V�4A��kK{��R!�E*�:��p/�D����"��(�$�j�2M�N���Lƙ��������l�{�0]�J���`��JC@��	�F����`����2�ˁ���]\j�k�'fC01��}�{[���QHE
-%�=s��^s�np�Ya��*�\x���W���P��J�M�B���;��t���~f�`j�Q�֑$!
����P������s?
�Hz�]#&����M���x#��P�~ �CҮ��C� �]S�ڧV��?��k%I�hD*��=���~;����V������}�B`��$ ���P�~ta�{��=�u�9���Ћ�³� a�����[!�a��:fY�X@?���"�G�|�r#	R��qʠC%�Wwy�����	�e����Q��"��I�*HQ��qe�i��s��*� ��7�9A���f��Bc�~|7��_�(��1|��k�*}(DܪeC�@���P1���>�֋Z���^{f�K"�ג]��TqCNLp,4�;�W=�.&lk�����}��N3%��EF����1� �`
I�Fy4�:��rIr,�&,�B��G.��	�f���XMAvX�����.1��Dh�(�J�ՠ�`8�TGq4�����b*��&�w�a˂��P3�Y��Ep�¢��V,)��P�:c>Nx�z�b*��UP�k[Wjp���3��$�ޛ/��Yl����xt�Н�4�tq	a��Ղ$�7����3^���U���j >��K/���C��l�0����*���;'�J柸Q_T�q��V�E
$�%�ؑ���Gj]'_CF����GIn陵��إ7�f��n��	C +!B�!"�V���i�@�)�^�$ٹ%���B�|�%��J��p+C��}̞�K��Q/0��{��Q���*`H�Oz�1��,���{]��y
#�S*����c	�Ze|��а)'���|e�F[;��Ĩ��y�S����o��1�;;�Ȥy[�I�0Q	I�m���ݺOV�]��.F�'�����Up�
��F]��7�US������EŰZ���E���-�ڰ[��ۋ��Qñ�@g�����f���ei��PS��;��L,����V6tIz:��ٯr������]i���q�����{Wr�g	��x�}b�As{M4�a q�c&���Kw���ڜ -b�ϐ��x}u���Q�����K��䵮j}x%}�Fh���Es�:��ʝ=zKM'v��-t*@BdkC�a���AA�d+G�����mWX�8����e��x�A�Kʁ�f ��#��XT�]�`���^qv|	���e�:�Q��TH���UvkWb�w;�c4yH���
"���t��t��_�ac�*�˅�2�٭��>�)7��ys��Ə��݅�`�#u�)�Ԯ-A�$4���?{zӱN����Z1��*��������aԷz+��T��p1��|`�9�8S�M�<�����U��S�,��Z_I���F�����q��Z"K��p��z	��uN�,DWq�epz3��r��9�}}�&��#�����u*/;3��ܢ�� �@9 ��$�#4�9��4���h[�Hn�/Y|S����L�_c�E���`��+�x�Jl��؀e�Hk"O+��h�e�c*x�j�xڐ4g��1�K�Ʉ�w�@�����#ZՋ�qgK��򈵁@il�gv> 	��bS�z��]ywY������:�=YG�8#|H'�g�>R*P�n��k%��F�-��
���!J{`q��ڧ7I�^s~	q�l�ibC��4���t�����S�{w�}q{񿢂�Io�<���5�u`L�B934'�Ȉn���{����	��GRR�S(F����y�;��Dy5i�U�,��t�$��tiƇ�M��t�ܙR��n���>Z!���'���ݼ�\��/�~ f({�����\��B����}�J���PS���*$ WMAe߻A9�~�LI23���Z^,F�Q�����7��C?߭�Vd�5FV�.v1G�6���T�^R�.?u��`�&�*���P��}�#	�/�1�o�f%^wb�AYm}:�jC�|�/`<� 3��
42�0|F�Z�Y�X�����&QG����V�]�'a�B�h+O�J榃8��X�����(�oZK�CΑa�.Щ��-H<�i���I�͞P�_�ڋ�Dǂ� �����(}�%dx��Dn���|#��\2Х���PU�h]G���HDM��y����K=+jA<�Z�zƩi-�9oe�	b=a@��+�ǝ��`�j�xl�}��|w>��F]+4� �|�A�6Y��/{ �팲�r�ծ��Ůl��F;V��1�N� 
=S�eִT;L�`˾2&�(�����x�l}��u�;�LL!��+���0YB�;M<q�ťׇ6u?o"�����(�C�������U��g�c$=oM��{ɸ5�T�;]I$�<��=3�k�Ӵ���"I�:w��������).%�_i~ń�Kxۍ�O�H^�#���������t�b�,��]Â� %����
�c�θ���C4��0º*����?�ɢ�o�'.����s����<��Eޫ�ZK=ԝ�Òĵn�9 l5�M��T��?���]��u1-����;%�����;��toq_#��O��U7���a
��F�e��y��R��Y��э+.��s�t�$�p�#�-��\�t^���yt����z�5�L��x�$��-~�m����Fa�k�J�0=��v�w	gUћu�*����׈	�#��X双��a�ϕ������k
@����}<sn]c{�:=�!o|fJ>hܤY�6 �2�K���/�8P���m}	eD�d��hM�{�Հ"�A}د��V@O{��&Z���0��aI�u7������!m��P���rO�r	M�����"�r�<�'v�'�"���P�Ԭ��H��6�Z���l��?�`�����z����������Ps�y���J��U�"�h0Y|���,�[�V/����M]����V}��.lojS;jK9����OВN���P��h�Y�{7�/&F���r���Ve=��T�]�����Y��Y����k.���d�6������W��:g���,�4V�_��`��3�3���3�R����FO$��j{7e��OK(��+�_�0�/�7���n1'\5�B���H;�Kd�Z	����5�Vn���j㚌��3
K��ǅ����輟�C:p�^�u��SO�v�X�(�6��^�Z��㌌�(��}b��y�����ҦV����,�
���5� �[��l9���/�[�L}��z���~� ���'�GXb;з=~��@��t�� ?��] ��|Oe�M���'*�t|�,��nw�D\�^��H�w[m��JN_�qsT�꘩M[\�@J����JpX)��������Eu�Z&�:�%�/`����h5$4�c��O����r�\� Ȓ;���^�/�3�x��`�De���"$%���kdX���M�Q8�y Ua&LM��q��d��6m+�����}	�O�_�����z��de�\�:�����Y�`�nL#�Zs�l�Ηv1�/�Z���ȪС�#7����z�Hz���ɱ��	����r�ѕg��ξ٘-�����AD~< ��D�t�6�ԗ(���2/���6������$q���p_�ђV/a�w��/)�����Z���m���B�����lϐ��#Tdҳ��8��l0u�t��T�\ֈ_�n깄{��sF�'F��� �:��3$��2��j`M|��{��S�����A2[��:���z�����%茮�������}���1j(-CA�hnt�ѕ�E���7���D4b��9�
dxV.=����L&ÛT�H�}R��n#�n[5�HЉ�cL�J��h���8|�?$z��9���<�@�=��z����u�c�H�l"k��ыja	
w��;��S�h<�'U�G.#�:��4 -o����{�P�Q�2��6�w�k	��3+�qq�!ǳ�h�
�J�Q=D��:3��II�̲�O#���˄�BE��O�p�n���hn_9�I����5<<pN�oec1v�o��Z��w�g���_�T����g��p��#Q���&4���E��כF8��_v��~ʷ���q�-&�C�pz�}�FGmFM;�V��ƭ���MӸ(9���͐Y�
`Vn�h�\[���4&�X�VD��t�2��LdR ���S���ߧ�r]�����0�r8�G���npd�J�7��i��kx�ɷ樬`:\o��cR��ەh(E�N�rO�.*dX��;��G6�����u-H�M�\c�]�.����*�1�Qá0��%m��U�C8���%�"�[��DGn:�ȳ�#j��>G4�cr
�,�z-�t�h�݁�Q��~����E��㻦�n����v��ҩ2��?�8];����� �vHԙ�oMvx՝pA�ܘK�uD��4����&������#dd������x�t�[�+�z�oQ��[�� �b����]������N���}g����VAT��@]�׼5�j�ڞ�sG�w9-�>b��f{>�z�z���$�b�S���9�eǏZ|0�yf���Lކb�k`��Ԋ��G����G��c��4E����T��Y\��sl4�M;�o�+O��� ���� L�ʎ��1�`v���ނ��(����Չ:��ߋ!��ٔ;d�98� e��C�X?�y�<��R���'�-2���P�(\��<���5��_=��0�uR��eh�nT�X�5��Di���G�Q"�ݼ����_/�5�uU
��gER���Q����CI��5�ů�F������,��6s��3N��u�}r��T�I~d�)��J� 
�L\]FNs\��睲|_5N��`}dK��k��D��2���Iih�e��I���I��Ш�l����S�у�5P)��(�X-���/�n��D���E[!|�q�(>r�����n�"��S�n}�6��N�%u��R��1@_��޿����\�ȯ~�نV^��[Kҟ)@�{L��lI0��|��2���sI�U�B_eJ�H�4�x�j!��ͤ<_�3+�t$LO�$�
�N����g"���� Ԩ���8�_�Up���1N����7DBD;�o��[9z�h0N�i9�o2Ϝl���O��-�$�*����h�C;|mN��(��w�M)�!�%�1X��E���X0�ɬ��\hfcIWǟ�M��*�v��΅z�.�gL��~�_	BĮ*!-����f������Vv�z � ]��������p|��;����Z���+�s�JG y���ݮ������>>���(��?����ɋ���I��P��	!=�I
)���Kt9uus��`lGB<��"��97t�������n´�����y���ES��'Wx����׼p�C	qSY�I��铛�\�u�_���eC�����bM}���y�s74>���ldU�J1�:�h6#�u�>�-@C�Uf�-s9��q,"��íA|�� �!����u�/0�k�#�n�ڷ�5�l�!֮��y6��=[Z9 ��9�h��xd��\V�e����\�$I�j���j�p�[�"��b7Jp��G�'hT��3Z3~L'�<���՘�Y�F'}dp94�$������$s�y\���5�߽�N���}�v�Ab�k�VN)����}���E�nX�u�@�0iaS��� �sA¸DX?���ok��$ڜ�@?pa�5����)�6�P��l��.ړի*�K�PK�G���Έ��I�^�K����Z��Ý������3c��NEE�
[s��4t�.�n�A���$�lf<>��_����'��6�V��I�:Lf�t��Y�Ym𭖋:Jyyz��&�q�˷A�(W�I"5�$2 i�[�
_�;l�7I��>&r�_��|��aF_���։$87EL$o���\�`���}��f�Dh/��/��ڈCzVx9��67-�{�?O/_��@.C`?�<!�\��mo��`�l�Čg�G�{�0��޸�B�S��m���:�|t��EL��Z��'�Ej�Ƀ4YoO���Ø����iaF����֊���s�aj5B`]C�o�]�Dze�U��2�R��,*[��{Q;4/!�brB
�6��j���3G�8Cv�e']ҷ����U!��p1�Fx�EL^�ɦ���C�̀�`�~��X�D���u��������7n����(�?�C9����V�Rݑ�=�&��Õ�1�|�g�W:��.A2���Ac�P�3i�$i������CHh�X��8b����P����X�~'ZZ�A
8+�k��26���筘�/�#.��U���<ֳ���YO.����8���;75O�|m%[Bu��-�#�Y-]�s�.B&�ߥ)�T�	W�!�1Tj���˃Qڝ����+�J�����>��J��g�K�	4����x~��S����F�|�8��d	?���i_�D���O~�"��O@)��5_H	%��^(R��-��%.� V��o��R�:��m4��%�o<@:�VR�~H����Kt�C���Z%�ב���$��؍��t��53!��g�c��1	ѹ~߫��7�~�}��c���D���x�C�d.vu����ۃ���D�z��iHEz:X	5|�6"{�&!ߒ�2g5Ф���������������݊
wd�cfl!G"�0���泓H'�H�X��k�d%
�U�bJ~X��nk�<���򺍟�Ǡ���A�o+��0T!o��4��?�/��tlsj��o�]h&��Ж��6:��jOEk����Y��D��^��Fk�br�"�=�W��	:����>Ȱ�uH����z��bBG߃�\�������f3�Y�+M��u�k��qB%��V��1t � +��m/�����G�f��V��-0<H�|*�0,��Zi�ᷪ�,�&��"W�TTa`B�W�a��'ٛ��$`)5��)(��+�H|O���]\�pG�%PѨ�c ^W��1:3�R�3.NDE����yKM崉ΧJԶ���I���4 +ӛMq�5�Ir~J�hF���Y��9����ԥԣ$~���j���]�����[����v�Fy�Ʋ�*��u;��Y�M$�&:��Y�������W�v4�@:f�J��P*��[���C3��zKT�w_+�Rq��ԲO9����k�L0�G�_�ᩤ[�I�7'`�-�Yl)MO����RT�H?g�u�{'ݣ/硚sسy+SUD��vm���g�YYe�@�]�Qew%V4%��\�.�W���-Cl^���s�(��b}Z0���i׬�]Z͓���p�a���	��ץ��U�m�''gۓ�8�~?�6�	4@v�g��v�Tu�<	���_+qH`Iέ5�9 ���F��g�V�M�S��.;vqT��{�;3��+QrL��b��c�@ف`6�fF�T���9�>(!<�B�:��^���a���}4�m;�e}���ȣ��:&�Oˇ-��4�k��\d������$*&#^',�'����Ĵ���b7aVإ�����#�{�kZ��Ng�K�@0!d�Ơn������S@�~|��W�r�@b�m4X�l'�([!�G@�jM���>�(�������8r�mu�q��>�w�\�Gc�4S{ҹ�P{�A�UHJ�����x�T��E��?�k)�F&�]���8a=`hi"wD�:�>K��a���׎��i���j�7x�:���Zy�%��
H�<�w���Auݚ�.'�6ԭh&�\zйыjK�G���Vp����=�tQM�ݿ\�릁`���w�s:Ǩ�|@l��$5��*�'�H'np㧏�W��
i��'T63�y�����B[�J]���2�@��j��L)�M���3�-sd[KA��8�
m'Ke�;�e+��$N�HW���獪-%���]<�ӖU���"����4�!����1aܽ�*J����mv+�a���1N�=���2�!l��t.�	�0V��Y(9��Z��ӧP��7m�瞝��e��T,xg���/��-m�a��"[��b&�����E����v1W����6om��ʹ=���d�۶�H�3�c�&���rrh��Q�V�[� �|,י��
	`�p�qrt�p�dHg�?}����_Qw�+��<�b��:���+�=o�`W�=��$���c="���s���C��2Z��S&��G�0�fQv(d)zf�����wpfq�>g��r^���BJ����US�4E��{��`���p��"�p�Б9ƴ�XVy�'[�Z:��ABrW鈫���Mm/�=�����S�/���"�؍t��Y�F��[�c���W���6̙�Ep�-��&�^��<0�K����w���	�K>^Ey�� z�m�珝�(
o�N/��d��{�~.E��;: ���/��ɔ�>VZY�7'%�(�J�NǛ6���QV/Ce�8���H]�p6]����}�g�h��:3��as�f2�X��M��Z�����/��ˎ5������f������d��$�$�)�PQ�����h�w�����jXXoR^TS|Š�Vx�	��P�Eu��V��=���y͠�L������/��"�w�M�UEb���r�mV���摺ā���<��h�(�Ʒê�����yo�,� �̸��o!�q�HgF��N�[���P��Cs��������JM��aA�%	h�M,˩Qdc���d<>H��
=����3���� rJL����б��~��!&:[S�S�^���Y�:qO�������=39�-i�EFdE>il�W��K��cU��q8��~�Y��k<j�_�u�ϖ
OZ�5gr���sb�m��#��H� ��
dI,� +��. �.Õ�[/��BQ��얲������0!�5 �(�+�)tza��>�ՎC��'�Hgő'ӘV����F7�۴B�h��f�,X���O3H]��o�T����NX���g�%�M�|���?�"_�D�+�E�,F����e�Ũ��^~���*[	D�A�su�9-D�b��ta컷`���{��Į��f�����!u���v����g�u�K���)���Y��vY�0��t.�Gb#����q�*E<W7a�l���3D Y��#K����4��=m巅d��[P���H�Ɍ�c;�fiHV��i1��W`�y�[�Z�A�k\�����k>�!���7�SǄ��޴��������<��-�s!��������a4
����d���B�0AGTH#�����r�(�9G�|�/'��t+��o�M�G�!�B�VC0��w����u���i�'���wwz�M�Ӟk�2-���'��[n�����x��?�\��m��gKݞP���������Q�r0�0���;�@H1"��_h����u���W`,lPj���tGH��SQ���BgJ�&Ĺ�p���~�|m+x�-��Ai%Xnnױ�Ɖ֏_t+�KK�doPjUM!ʛ>���D�ǹ�ae\�NC�e�d?�7*�Hi�x���7�24�RF�d��m�HN,�O����Zג��
�%M��<A��%��n� 
�p�d���u)g��B	`���b������t���OuS��WDv��$I�*��0x2`�}b�$�D�j�GDl〣�z�ZnC�N�'�>g���-
�C:��,h��z"Z+~�<�%\���ǲ�,%3�������rc1���`���(��$#�1�n)3��3$k(�v{����cT�@BZ~���s��^���ǳ�"�� Ƚ!1]g).��Yss��LG�r?Uj7��a�=VCH�����C"���ko�4q������R�'l⌖r�v� 8L08��/&љ��DU���ƿ������7��?��>h\7�K\lb��� �S�
���&K���^1l�/䌡��O_;0Ȋ��Я�X�`lJ4��y�?;��^e2jxS��%ꀂh�N���s�l���z�2��vJÅa�����=D�|=wV��&��܎� ��L ��.�����-a�*I�Z�ʬT����9�f�%�>��!%|r�ʇj�@�Pj����#�U`e2�́�Rg�R�ups�f��Z�W����3�0�*x���GiCN�n�*�n^д'A�z(ҙ��@=�K3rԒ`�h=�6.�y嚿s���4�\;�#�2&�t�q����ko�1ڥ�{7��X������T��K-��Ǟ����6�T�"���xi�;R�}v�f���^�>�mV��k=�IGŹ��rs�����D�����������yE�+Y�[�yRMD�5sʆ{Q��e P�|���p�ѷx$ ']s���c�E� �}���s��g����mƑP���ɆA˯]��;G͡+(U��&1�'G���2�˨O0_����[K���9�M`�ɦ�ui���^e�c=�������"7/Mo#����Hܘ�=x��O��	ŉZ�3����$��?W�.:�=��-����3���sw�Kg��$�w��be�&��2�5���K%���H�#I�0R߳D���5d!fDų��	,][�YQ�/P[o�oZ��E�Hi���Kn>`0�4�ȏ3�] �lz��<��<Ƴ�b�3�/��[e���(X;�pe�)C�"�s��g.*r�z�+��Y��<
	��E?aJ��>��'�y��c�Gto�}8�ܫР����D��z�ٝ^��z��$��5��`)��݇,#�T����m�I��3����U�B��4�^�'K�吗�lQ���	6��q����j��}|���꫆g�f{����n��H���?1�{�M��F7���*M�*~�ǩ���tk���[������2�5�B)�3�����q����X���;yU���j{s⍪�mQ��gT��CY1��+_q/�hJ1�n����8�B gӳ}L<*㵡�D�"1�^;S#_(>�^��b�{P�oJ��yZ���P���|0n�*�2M�Q�t���]@�HI��"��ġ�d0��ˎ9�a����k�G#7*cX������k��$m����5T:�Q��h����HT#�����̵�˹�q�6Oq�6��&I���|<DE�����b�4r��]�A�i������kz:��6�B������`ɿ��ﴗ��*.�.f�|�pgQ�#c;�\��N�c.],��2�@x5X����LF��|�LD�ý�:��9i9����O���#���;;�!ƹ	.Զ w\R��_���Gx�1�b��`t�M��V�C��������%��Ik=����N�A�=62_�ݩ�'�\J�<��H���!�J�8n������n
ҚeO��`raz��+Ρb�7% 2��P��z���`o�)ai�y�h�>��q
=������v���xwo���q=�-�{�?O�� ���8�(p��#Ֆ��Vf������m� Y�V6����x�� �b��������u�z+ʊU����ɒ�����#=I���<�V�f '��o���N#��7p�p���7k�xBZN���M�dѱˤ;��M�\�> ~�4I/�W�gW�蘼���z�~��$�p�;�(��⑊7Ak{�9e^��)Y��R�.FU�ʺ�٪F�u�J˩sA���J"}�W1O/P�L�������p��]up�Xo��²�'�-4*��[�b���0hY+���b�ͨ�D�G��ɤ$_E���/*�v	��
��Oet�c6������?F)n���D4�,}zPج�D��痟<��{�K�a���6�؝6�pN����';�K�d�1�������+�[2��S��`����!�X*�>HsTP�_�n�4n6�s?��.*���Qe>�W��/蹮�=�NC�gy�(�����'�����(�i���(�̫c#io2��3���h��0����W؛R����Qx�EX�\���Xd����l$/	�]a*"("z�9�%��%<=�S��s���&\'�CN�{�܈H��ê�WΕ�uo���_I���;���%�����ĶU\����c��zL�GP��J6���|��u� �8 �F�窵�e�Hs�	�ԧ�A�ј�Hg�����M�ҭ�ی	�s��K~�q�{@����jA��_��P���A���:�g"2r�-J@<�����N�,��_e�-�&C��]F�q}�l O�C�K��N����U���<���i����lo���{HD�����;�ݶ���K�5TS=�0�N���Ϩ��D/����w�3v��,<�b�4ӧ�$��˾?c�v�P� w}t��Ͻ�T|fװ�u(W��L!���a�v�/�<T�h�ǒY���d'{�S�[uW��>��b����}��A�� 
V���9Z���)��ou���]�p� V0�2|�my�ӥ~��=+���n��SER�����G����W`kqO[��V��9���W뽼��aq�`�7�f�-�a�T��QE>̨�~M�ӳ�+*��Y��Pe�����������3G��ƖZ.&��$� Us��Л�	��|�;l� �����LC|�!gq[&)���Z�.K+�.�
#C��T���z�Wy��_�Z�����;9��A!:�:��c{h@Z�o��]�(U?*0�����{aI|���!�}}���,aF{`|�����1t��<��*�m7�ھa-E�8���ә��p������s�x��զ8��@)��B=4�;N����I���~�`�HW���]u�����z}���3H"|o�I��jh�:ؖ���Bb�\c����~di���dg�s!�a�>��6cd0����T_bf��g��oKT`nDD���+HG�����ߦ���l��-��z�e/D|��6*��C>��ʣ�R��涑z�G��T;8����Fģ*$C+�᣻G���Ҵ�FV̏'?K\2i�4oJ�"�e*����l�=������Y��с���=x]ax�T@��L�7/� =3@�Mvj��� h$P,��W@SB�h���Oȩ����x��1�3���o�5�=�y�Uh'��f��B�3X�.��f{L��w����B�&=�`�b��2�����Fj^��v��k@?g4����zt]y	֎��|��WJI�Ck����X�:@�����w��g�-	|����L;�4:�d��l�cUA�9?�B[S2�Y���;��Ʀ�{߁%t^_^��N+D�����#2a�4��[tt�5wTCc���s@<W>�u���V��x#����!]CK�ϲ:W�M3-.>�Ң���0�L���ϴ!Y��<tA�,��kfeH#p�M_��4�O�:E�!��"r�D�,M���&�X��s�@���j,�k�O���Ǡ����A�a$��g�Qc��d�dh�	�\�]�I9PP^�'�6V㭿����#�­�v�Kjb���կA(G�*�g�����l�c!��ȢMYL�y�pe�����r������p��i�12m�޽�c�#6����6Z�>2������Ȉ^J��~W"���7��#o����oÉ8wZ켢lDE�������N��OH@FL�NmV�� Cw�=
����Ƿw����0��dB����?�f�����1�LB���3�ݚ�_ �����������%�mc�Z�Y+\�髿���+�
�pz26B��25����" 	�K�#��:I[�f�_T�n���8fۇ��g"�bע?~��#<:�q�R�bS�23�g*�WxX�*	�/�������[����0;ղ�����S�_�f�f����t�F���b�N��Y���p��wi�Vq�>v�iT>��R z"g�6&���D����U13_��H�*}h�(5Z���L�_�o�s��u%�}N�w��7���D���N����&�H���:{�T��u�}��:�Q��̐�v�+
�(s2��"��l�.O��J;\��H�4����+�RQ�@���Ȩ�QCF��̨4s����A�a�M5ڜH������UJ��!o+!�Aa,m+�����!)�l�!#�Eљ���q�)L
۞k���q�[�GU�B��ꏋW tȂ`�ٽ1qZ
)��K*lAHR�U�K�֔�j`�-?o|��:�iT��Yӆ}�x�}�����Ԇ�ⵆ����2ZC>o�E7�v�L]���3�81+q�Bڏ��=���
���~r���}���l�k֭=��B��m��Y��R�����u7�#�n�
�tn��P�/j�X�+�m����@$ר`�TC��F����JQ:C{M��+�Qg�r�!Y�N5�=`���	s3��]�g�)B%�XE��ii�1��q�*�R�Pvs�9�G@;�9�b�1�A&pT�G,�1�$Oi:OBV$w�tD/�n"�L��x�%=a�2 4���Q�?�(�V��}c/� [���W�#.!Ã�i�2
;�YmֱMyl���H?���ܦ�d���/�! ���P����s�_v���s5��Ǌ���W<���X���ʠM��KO�W��HA��R`.�yv�]���گtl-�����D+C�*Ԯf���F3�@��G���*���F���:a�R�>T��`��@�����SX�3�6U_����;����������yU�ˏ�(�C��26ΰ�O�����D�en���g�l/���v�v����m|����ry?9��D�A��P�ET�W
ҡPK'VX@5+.���0�ӊ��{4!m�� �m����9�����x|�l�a�NKP���m�t�V�U��`#�V����2��ί�#���x>{�샺��� �<7�����t�`G��3�N�Gj��t�WU��/t��� 1_a�R�\q���k��5�;fa���x�Ye���m3���{.�;�f�����1��<�z:ʨ,ɦ�Q[`�N�G��D�� wa��-p����`�D����� ����@d/T��J�(�x�I��'%6���B���ԤF��de��re��&��C#�uN��k��3�R��lVc�e���-��)*�p�2`�-z�%��/ě�{�8MG���J凁u&V��z0���>���������Ip(q(j*�v ��5�s�nYo�����|ģ���5�	%�S,|�1^�SV	��rF�D3Qf��sU	�#0 `�jR�t�c9���TQ��%);@f�F_��wO��6�C�h�Q����ø��X�V������P�U��[B	�{w!�i`ǐz���Z54��6���&̍<�Fz���E	���uăg=�n-J3|g3��	"(��A8�Z���<i�����	�h߲ʹϞ�c')X
_!+"9�ǉ'�����`8���PB��L�c�v��}ʗ!���*���Eₜ�k�cy��9�پ�ã�Hڧ��ԈͶQ�x0+���.�G�bŉg\Ka�ҏ���7� (u�d��\�����s�:ݯ�W���!2X�&�4>�0R��� H�e�C&7���Ӗ&j* �4R���df��/�|dU�b�`@���{���y�
4�Xd�9�N��Ʃ &��M��կ�wh)<�qۧ:Gb��eϊ�0hm��6�����9�yf9>ߺi,��:�$���K
&�}7?�D��}�W�s��5��U{(�T!#��ŀ�܌DX���9� ){C󓌕�9g���e"e[m����o�snT?���J�\۰�6EW���j�3�͎@�{Ӯ�����Ȍ.�
�#]Q~?�i���"����1���Vķ!�]�,��˨���{�r������\n̕mEi���\�����W���M�gc<���mS�ûc��Zw����8�7�R�?~��f��D�]CP0�x����Z�^/%4*�y
�Q7\a �eh��o�W�Jc3R�[��fd�	���i��I:��C�
<��q�Ӂ�;ʆ >M 9;���B��ޒ�lWu���v��O�����ͦ@%����j�N_��f��v�{��퓬w^�z��	I��m(�fu;�E��oo&�֜ ��(�T��uĻ�����D�������%V�4+KH^��vgG�k��=$�a�?4Z��E�M�ڙЕ2�.�����~@ƁIGgFI,v~r�y"?�����)����t
aMu�súo��D�=8��r�a���ǿ_�fk��� ��Vɵ�URp�-�T��ٟ�|�(1.����N��]�HΑ\]klx��=y�g���X⸞���d��1RR��5t+��o���y^E=34��܈|m�$����}h���g�x��j�MF9�Ț#�a6�r���h�A�ہκ[0�������\�qz���oS�1��ˮf��Fd~��/�&榹
����U��m4���A�-_���/�}0�E��ľA�y��c��Ӷ,�J�4�����%�..��j1	�á<7�EH���f�Nk��Z�Q9�4//�B�B��i=���h�YC������u9�{F�ܭi�Tѕ��^�f���#
�F����q����-L���=9,6�o��1��P����lN0�21�\��<eRw{vX�}=��'+��Z�F�.Jւp�Q�����
�B���0|�Gq&�8gy�����$����W?�]�%��cwnUh1m!bI������'V���X㛝�M�2}�0@��3�U	�|�!��{[����X%暛]x.��^�w��0,����پ�~�Ԩ`�%e���
�L�h�7���[�T��Ԙ��ɀ� C:6��}��9� �`I����Z}�Yqw��Oۏީ�?�R�Մt)�a����3����X�u�`!�+nqP�#�+WYLK��k$��|F�W�+ڏ��� )�
zk��P�-�Pָe)�yeOܓ�7�RD�;]�Y�Uy2SuU09�1ɕ�omY��u'��gz���h��Ja��QM#�y�Q+�����
&��L!}Bٱ�6T�F"`,�񍉸�.���@�u|��-���j��/�)^�����ܢ�J�O�I'�ϷW�PM�華�_S?�Э�\'�?�9l���.�|��%Z@�C˯D��+�]�����w�|Dr#�-;ۏ���:�}�����݆�<���ǖ��Nթq�,�m!|ݭ@FV�IPØ��,_Hw��쇬�qg���H�^_���F�k����`�+=<s��v�vm��y�`悑n�\�"V0�h�wtg˿���b�f�d���u��ݖ jJl���g�� ���<�G��B�떷H~
�*��$�7��?,��2�Z>��a��|(�I�N�*)�}�w�@.�?p��I��AG���f�Nb���ޒ�,\�w�pT�̈�]�O!�Rkq���z��j�,[bVO�!e��q�b]�s�P�o[�
Oى?A��AhR��,�y7�f+�Ӯ2�D�_Rg��ߗ�~��`�o�D���.�M��*)�o�Œ�s�=��v=�)#���ɷ��˂�YD�J�	���0�P���x��m�<��$�<���W>o��
vQ�ƴx�ҭI-4�&�,�P�����*�ǩեY����} I#������G*i��W���@�D�Η�j+�GI[�L���U2��_c�83���",�5�mzϱ�d�d�-;Ѷ����ܒ~�q�Z�p�87�/$���2 A��^6���]�����=��W��)Dz��Y�\�W��O�xތ�;W���ƕ�ͬ
E��Ѳ�C�J7��Zd�i<Ǐ����'�f�7>Z�k��o��뮅8+��-"�굌=C�������7i��n���Q����#I�ѩ8����tN���L�$�QB{�	�����n����UFɘ!�X��.�l5��%(&��3K]� 	Ƀ�����D �e]��;cdq��D�vn�Z>6�H�����i���)q:�$�ۍ`����8�Z#��E����UIc��핖A��U���m�*���G6z����//�U��ҷ� ���E��D�feV�z�b��vZ3�~A�r~��x�6������U�ߢ,���x���X?�������?�kk9�H� ?EG������HtS2��� �z�j�����y\��I �G��%�[}��nD���WSGT�,G�g�u
��E{��|�%�"�w�2�&�@�'���c���(�D�٣�������΅��GkJ���!���˃��] �"�6[$8�Vՠ�|�`�Fg���'@؇ڦ;�4щ�	dy@��Cߞ�w֐����<�g��+�:~�t�g��{�en��y�8f�� KK��|-�P@�6l��jC;_~8�O�b��r�HYI���3K��d�k��»�� ��5�tl���9>�Z����Mx� ~�xY`��J���P�W��q缇��v�����"!��M�����E�v�u��wQߨ��Ͳ/ډ��V���w>��GH+����^�0`ZQ�\=��<�Tch.�A��bnl*��1{���"���.e}'�ZO%�I��T��xS��S ְ��욬�aGmj���i��Y�i�S�/�� 4�p�ɒ�I2�,�
ٹ�?I
TNcc�VߏҲo�d���V-�jߕ ��H��B��Sz�w��l�iĵqoK�n6
�K�-B�
'�\��+�+_��Al�'��i&���Y�����U��J9��p�(H��T�i�Ȯ"|��� hΧkG{1ጪ0�����Ҫ+��tA�Cb ��>�����Q�[������p��CE���%A��8%����W!�Z��>.�\[��+A!vj,��@;��A��lߟ�0�~f8�0�!8v1�'y^b#aA��q_�y��*��v����F�˻S��T+[���JF��J�_���L��2[0z:@���J�,K7� ����+=ӣ��xA�<�1޹�S���#��ev��:��L�ȶ���5{�)z��2.>������(G:�ou�L��3���d3���D|A��c�i���5�|I�	Wk1�h�5�K���'Ai�����0�G���S�3.�j��]��`@�XLy�'���{"���yDmE^���'n]=��.&���=��
���p�j뙟/����~�SHU�	��*�g��#��_�c��q�����#y��ٌ:��Ȯ�� sj9��wu{��䝲9eI�e�4����������=7F��T�< !2?>�~sn'�59�ul���b����u>[��O���4(���PӖ�[�)O���H���z�����wW�Y�UH�2f���d�;��*�!h�l�ݻ!"G3�^�Q��Χ�f!؀���]���
��)(����4g����=:;�p�
���#@0��C��Y*�F��O��i���In �6�&�ק==�kL�;��}m���q�Y<��r���y(� ��\��)b���s���q,D���j������l�i �}��W��Ċ�@C
q-�OSW�u�t,���ȋ��ӣRaxe��A>��ܫ��� =��5I�^}�0�~�$=�ۊ� �������[սU��
B;�5��3H��/������--�7��p5;e��V��8�&p���"�w�3�Z`����6R�Q�%�ՔM�z+�r��Z���D�9������{��X,=����t��e��϶B}�P�VF�{��Ɩ$3{\�F�KbΈ��X>ud�,7 qEI��?IK)A5ϲ�6�fuV�ȚJ&J���Z`�E�U7�<p�LY�鍂Md�h:p|y��7���	�.�����Ff�7������:�I��Vq4�Q�J#�0�TV5O��	���0����y�Y�I���g16ˆ:A�un<}�}�_���$4Te���!�����k3�3�]+�)��?�2y 	G�ڛ��z-O�Zu�D�'&�{�����I逃��z���T�>\�k���e PZG�/����/�Ч�Ӟk�|��hq=J�IP}9(���H�E�7�2�u�(#�N�?���K��W,bk�
ˀ���kF|�J��W�v(�A ��<�uѪ�K�����{��]}zԝ�a��<��2�1?�d2�����Ơ�UA�������J<XAB?2n�.������y�#K�����w`���/c�,�;�W���T)�[ld��-�Aɲ}�9�mP����j+�y�Z㋴&Ŝ.f��-�+)�fo��´u��=�N�݌���{��S%�7�6���A&�T0�X"��!�IIZca�5�E���[;�4�h�?wT��ߓ\\\�bv���vO�s�����WѰ%�w�]��>��f�4����
/�\"�L�&}ժ��8,�c8l�T�w܃��$���tp�ɦT�:d������R��h��=-Ȅ�%�ы�y �������%��n!i�>�}r��1Dm��h�i���9��\�B�;+��Geݤ�`6��I5�X
��H���Ac�lJ���m����b���K"=� N�=5�i)�{R(���#�`��X���R�N��2]y?G|��T]aW'y�Ξ�;+��+�#s�;Y�.`%[�_$E�r@�����WIdz륇��3N�b]I �n@��ж��i(.[��@�+���{v�!��CP�C�V s�\����l�4L:�K}�O��߮5�{�����[�o�t��fiK^��R�B*�>�����m5�@p�1@!���T`�G���-O�RȜ�k2�����w����4R#�\��V����r�N� �>cv���/aV��ȏ�/Z���������_��1cL���L{���I#I,�8Bs�Q���$��A��*;����|� 5n5^�a<+�C�k�L4}	�z;��>��� E��F�GM� ��$����U�v��aN�D��;���k��w��2u{��2�� �����2ynҗ��ƞ��\�O(�ܝ��IBZ�_�T�z�f)�AJu�C{ǌ���2��p+�^Z���\L_g�2�����,��,XMy�B���j��+�-�Hwh�*E�B�"%��I?"�ub	)=h3L���yIR	b�HO����`qJouTS'r��k��==fo��G4��"�0�h�����ͥn��Z������?
kFh��l��Gw=UD+3���'�90�����*�j7���Z��k�ն�KFs�U����n ��sN��u�{3V��M�((�Y/��;���K29-3���K[���غ)e}�":�O���C@�[qԊ�~�-��y[*U�ug<�VW����KA����c�����~�ߣ�i����p4"�BYKyN�ɾ%�8(֯�ΤY3�"x�z�1O�P��sg�2�O^`���Q�^�������/�<	������æߡ�:�*g�yE��*�G)�Su!�rM�ȧU�X�	*b�!9u�wz�ݹyC8���H��	��a7�ZK
Z�6\�.��glgE�G��@�=��o�8��@����a�D�X���_e��ڄ�΁cW�)��[��/�=~F�U�MJ�N��9&�Y��l��__l�㓙˲0�taН:f�;|VJ�t,�G�ת�m�#}�|i��^���>��R�`a�����[Z)V)��P�5��_���_{���D`K���t�zh6z�,AJ�@�:�|�e��'2����+�;>�r�'^��U�c���!j���m��0��[�j��{�U�bʈ��;�)����f��sS�HX�I״��~3L�< ��>[��@�v`]�]f��w�I���a��(�]�c�)�~������.,@�p~��PU�����X=�/@#3e���뇆�WJc��y�IN"x{���,�X/F���O�Jgݏ�������f���jy�+_TQ3���twI`�A �log�&�鴡9&�͌dg0[#T�3��f柁"w��pB?��u|�VL-���QN�M+��J�?�v�P �}�GmǏO�>B6j�I�T�)ʫCx���?[��W�֪s:�RH�Y$�Z��●�Z�I����Y�L��n��
��뙍����êW����tk�����^�άl�v_�|�L���b��[������6){�I
y��x�<+w��AbI���^h�['N sSRٚ�}����95��*>�{v�2&[S��;WH����� �9'i�A�*w��/V5��R�i)"�M�ڑ����9�~c���h�*h�=�K.���̦�q}�"���5=�A���'�~R�59��]L;-.^_�ՖFGX�K0*��¸4`i޵Sm�� � m�Yz��G_N���C�_{�
F���)�
��h`(%�'X����O�t$KMpq\!�-�R�������+κ~���M|�ጷ�5��t׹�H��r�1d��U��;�ֵxz����G�����j!�y�}�0���o62�������Yh^���ߦ��������"�VJ��JQ��O���}x�u����4~ ��=����;:\���$��CN����[�!�5�7t���{O��()������� %#�m��-����C���-(�@_$bf�暌���4�mp�?�} .S�#SL�m�\{��Z�6�y{��p�)��Ѭ�J0J5+Pi\��f� ��g�Ç����5b7�Z�yH�s���+
NyW�cGXQr���V���qn7������Ò�ۨ����+��b����,G������QJ���t���Sm�����S�à+:��͢``����ȕV{s�ǻ	t�w�KIA��^Z�fz	�	qr�	���� Uq�Y�7�/�I�3�������Z�%Sn �kQ�A�u�aJ	2�{т��)K�TvB�?Ir������,�OX+�/�y����Ir��w�t7͝J�F3Ȧ#Q��?,��/R�`���.�����Z�H�����=�.��SGR�6[Z]U�/�>g����#��(2�0�U��q��m�����*�e?�,e����	v��$�t������^&>�r��`�����xg�| ��3Bǈ��M>�%K������&ma���J�o��������57�@6̈�P��*��2�5K</�-Dխ��?4���Z}Ғ���-ǒ�\�q��akO������V��t����	2�ף��,�4"���kQ�-�j���oN�3����|�N�ů�0mo��0w]�{�<'HE����Xщ �W�	y~�Wo*x�"�V6+T�����~�M[�Y�����ͻq\�EZi�^W���@����D¥(�ֱP��:׃l�]93_��ޖc�V${ޥ-���Ĉ��P���3t�g;�� ~b�boP b9>�*�Ǘ�.�9���hC�IN!6L�&R����#�
��1w8�+Y�q�������J[���N3z�#�@g΄����b����ضL#=-�'t��I睅a�C5��'�����؃3k�0e�/��S��9������&�йXnݠ�v
�����$/H1Ô,+��&��{������2[�͠�6O	HG���Jp���]e�����)���Z	��@ ��Dĉa�y킐����R���e'��kN: ���Ep2��[L�dS�+�@������B�u+/�f�$�?P��w�@$�1�q���bV:j��u o�\��$|i7��.��Uȸ�n�=��������%	C�y��;��zOf�����m��h�+7G����Cԋ�j~؛�۾��K�t��Yz��%��"Sx�*��W��ȿ9��%��̯fx�+�X�OT�%ܢ/��.w�d�1m!]������W,��9M�1+�-�TD���7}��f�>�n�ם�-��e1�hhE��OHȋ�E9T_����'�2���5��
�Wҫ3�Ʉ�J�	c�A�=Օ�6�-�Ҝ���L(�W����hxiм��{/��fX��ev@I3ɳ3)맭���Ν��#��;�L^�H/	����ѣj����e���>&���
������#�T��f��g�b����#��ӆ�KL&����e�X���G�$/R�%)��NuC���^��ZG�XA����[�� 0y<��B5���"��<�X���ꋧ d�">hI��>0�;��[��pN9��\�o�,
��?�D��g��x��.�}��)T�5v���m���g�;<�K*�7�¸*H��4k���!٭��c�t?~!�P5W�҉�:������\��1�M�h�YQ�X<C�=��q�%&S5$�����	�O�pzt)�2�OH�Ѐ��� |SD_����o�D�l�`	*�������K�� K�Ej���T�g��>Ԩ(Z���CD"d�f,�S����k���{���b��g<�Ir\��P#�v0��� �����Q�,�W��8:L�ÇR� ���Qõ�����>FV-+.>���m���w�]��f�|KJ�r�ݻo�	0��$<�&�x�Cw��0�yv��������\&b����WO��{�Wq �)�~
qT`�����;�����G} �~�%-t�Թ�LW�C�ub�m���"���p�8nbJS�r\�T���������
8�I��+wGk6����J��Pa3�B�,L��I�F�`�R@:V���%5�'�PA�?���`#����P�>g5�sxW%����g�sxt��X���ΰ�a���	t ��k���İ ��}�I�����;ebi�h����Ư��0f{��|;\; �(��.	@a����uE��3�l����H�A=l|h�,w���?\�	��Vs��,;5��AJs+T���0>(��p�$=�Q���V�Klz��l�~�:�%p?<�yR�xЫ��+��@%��X��>�n����C$��X�6�ň�UHM_Ǟܞin��,݈�i0w�t�g���#5���T�'���B*��O��}�g9����!���G*y
ۻ���͆	�Snz� m��q�ٵY�֮o��o�*�������7ƁO��G5�(I�����P���&1o�,�ț���9�T�1��$I�����s��CW0�ㅫ�Dֽ�(�t���p{N���ү=���ۑ8"\6˭.{G�O�y�����D�� �T�M�;7}��q�)Qyq������e:o�ш�9��T�?��oD����.Y�]o)̩����]W ������i�r0+x�v��EE�î��b_����I��e�k�dҒhe���k8+"`��,�s��W�<��R��M�BBfg������¥d���ԝ�<�:Cm���.`3%5��������oG�	AI�B%�*���˧�ԲV�Y����������F-u��F�6춴#h�	���D�/q4�?����6���=�)��Jɥ�
>�� ��M�3y���He�K�f7z��������@U��,��z��B��ޠ?���2�`�VƎ�����ɔW0��(-�J��y��n_ZDV?��Jg���l�$z?��6�XS�v�aB��et6	�{�S�^?1H�W�q�����Vk���n�J�Z��h� ������;r�vfQ�9E&�2��픴���Y�,:�a�FP�}ɇ�p&ƺ��Y�����O��e1�N��U�@fsoA���ss�`�]_����&o}<�P̸T�8��!�1�p(Р�Ԇ$�o�KҎ������iz2EԈt�t��Y�,f�>�#�!wK�$��P���ju����~������/��h!�o�ʷEx��Z
!���Lq�Z@	����
�2�C����{��ҳ4�<��u�8~�����t��o[�5/���1⤮���Y�&���rAd��ݚζo�8��v5x���7�������bQ�^��_��m������
���q�qY���k����0�]��T{�t^W�錉\��������1���S�x_f�k���4����҄���1���;a�G�c�Uu����sD����I��N�MU$�0�4/�g�pß�L��q�D܌>�.����� j�^2�� �'�4�Q7oT�VB��ʺ��Q��E��\%�x#���b!��G"�n��l��Q7�	n%�[e.��#�Fu&0�r�*^�jk�[>NsH��4�Hn���cPm�c���r#z�O�@��P+l{�<:��;n�zc�F,ar_�ӉD�d���* S��%mbC\��ލ0>��PBdU��Ak�ͮ:��V0<x0(솏>�^�y��=�,�F�b���++��ڛs&���;��dV�K��,HsE��9�������աD*+�N-��&��*�	�&��H$�����4J]LcM�A/�sXb��z^�����a�s�������{�b��k�=eد���ͫ���s���HT��~)�o��d�H�ĝC�:�iqu����1�5L)��gN��7ٶ�r03������ �0���$:�PT���E8���u�����t��`�5�3�b�S�T����B��2�	X���}��Nw��$�nQK���x��DO�}�[�r�� �o@��
�3~�(��_^��������: ��%�S][�w�NTR�Lz��wi#��X�d��\���
�a�J���p��rt��̑�L�*ߞ��[6<��^r[XeI���ci�P��ɺ�5{{����?(
F"�>N[A�]���0��0'��C��A_��B����,�ɑ���q�j��ݸ@���ӑKr'η|��(+�D5{1c)F��m����r*�)������X�Ĵ��[h�Y�i�&>��ϑ���;5��Đ�f~M�>�>��Չ(�#��`��nkڬ쀠Uu��(��ᰒ\��J��7�Mѫ>O���Zm�pB:a)a`�Ԁw��Uc��3ׯ����ڳN���A?�Q�h�� �H�&3��4(�2�Ze��Li�ֳ���;��e)���A�׍��e�?���%#�CPȝh���$7^%֎KL�N�TS�i(�`�j�Zdcq�Aҧg�H=,�b �K���+�d�|�k������������d+rɗ��9RF�.�X�Tҫ.Z�U6ab;�������g��Zo�m�G��Cm��Bʾf�><C��h
yw2�"�3H�)IdG��Dkf�'8|�A�g���9\ ����ŖLI�Z��*��i�E��N3����L����6]%��@O�� �^/h�@R�A��y�^$�a�[3�O�!���F4���:��(Yv�v ���+�4ヤ�)��7/#g���!�������Ũ�&��z!�Ғl��e䘇\�1��'�/�/�͵Z�:�r�Aת�@�kf�FL�\6bX��fU+LbҲ	�S��_��z
k�tS&�Ig�6��~t7�ɆO�%� ��/]�:M���-P��j���硉h���\,]~z�S�R6���gD�,�w�U����
3$~(���^z���e�k��|�ihC0�Y�?XC����rjZ"�� t���.Qb |�1*oܣ~����-�~&z�FC�W�d�"6ZD���g�:+���R
OH�ʼXpӑ��J����+�HCM�R�a��6�N9�XuZV:��*�#3��7���u��&O6D�GrF���
 �L��O'�G{�Sk����'�ūU���1|O]��b6h6�<al!�y��$A|NY��J���� U���6Ԗ��ZĻ�Sw���T�C�WP 
�Z�d*��fe��ǩH��2X��
�	�K�|�\j(����~�c-�T'6�2G<{R�"�(�����-~;ђ����?��b� ��T1��N�z�\݃b���:�A#�#���wy� a��R[�B�Jxؓú�S�R�n�ӆ@���,�v>[�lG����(ft�����2����J��Y�Q����ݲ޾�̈v5@��e(��a<Ex�5�����¸�i�ܑ� �$�s��AC��M�с�#y�uMBa���3%i�%O��Ϙ���Cq7���>�^��^$����_4�8[��5"�qPwh�`φ�����2��������%E]�ǭ)��T(Ӽ��N���j�����53�$4a�0,�D��H�V��b��c�ݩV�O�9J����	� �����ǲD�j�?^�Ŭ�%�Q
� ��W`gz5�f�y;_7��F�2;٤�Xei�� FZ�IU�{W��	M��Ў�~/"yL�&�P�Y윍}�Ki߅\���91�;��/m�M^s�7nd�<�҆�N�����u��l���2$Hg����d�T�鲌���=:���t�ÅE�1���9Z�X��@����撿A�ų�=�J*�X���J0���Ȭ��J�>z�P
��ïua��$�2�@���c�	V>�K�im��%	\z���QB��@�����Rv���9�٣r�<0���!lw�[�o�g��H�W�81�33��x�VF�Q
�RCW6ۋ,�
��y���w#���Þ�rs>+C� qw�� �A�更T����HvrU`��ź'�� ���H��ȍ� ���FN�!����0��%}��Q��K�r����0i/���J�n���;��]��;���c�L��5�&U��oj��Es˔�|�᫂��u���=�	)s��f���6�x�ٹ��Cǻc�Y�D��Ő�(�B��i讪E9k2o<��EB�5Q���h����_r�vӑ�~��	��&��眚`���20e���&�������]��������̖�f]���y�xV���'W����1�S"� ����
W'�M:��JrS�p�E�<[���Ѐ�\	��'Z�ه�vFHc:+�Y+��T��Fވ��P��k=��c�|� r}~.�@��{t;�m|��M���DY4S�l��۬<p��nr�j+ڍ\����2�"��'�y����MAo؈�`��Am�l/#�(�fD�!tI�^C0�y��&���	���άw3�`�����{�ݰ�S� �254���e\̎r��q4h&;���7���s��3�bG�k�73��۬+,�Yɚf����$�"����iӂbGIW�{���.��{Bq����9z�q7\��D>�n��
��M��p��#%������W��H�߈6!<��U�^�,Pl�9�*t+0��8O=��A<ۿe��P$���R;�3fH#��K\'}m��5��f�������TD&�n⯲�sH��Y䫚 -}{3����KD؄]����/���f��L��`�k�^"���X��ܐ!c�����>��3�G��W3>)	(AU�_@0��g�3N�n�!�*��=Ii&>��q���+�J[=�
�;���<ef'%��PV�+�<�aq6�z���t�5��|�|��K1+�⣧��R\ּ�)�>�/"P:fv_~U��:��OmߡBg���0U�b}�I���m|���J�GD�m��	���X�݅����h��	Qv̍���A���d��aG:P'�����b�%���x�}o���:!�+�} 1��%������	��/?{�6hu��\���g�<V.SAf+Sf�b9%d���.(m�!lY����I2y�|�2�o�U�Ѫ�B�A�W�xXŸ>N/�6�'>jh���n�)�� ���V�%��Հ?�B$_�`����}c�!��R���GdV0����U�k�
W��d��/]���m�Eb�(�E�v�FYzm0�ɕ�o��rD�_^%f�P_P0�E����H�����!lh^�$�ꇹ�r�EK�$����}|�]��׌o���Q�	�X�Z�Q|nvq���j0c�}��5L����Y��ʝ��\Nw�n��xnnC�W�k��r�{(�}"
�����D���:�@B�8�O�|C������b�'��d�HaŬ��4�y�ҥă!�Җh��+E��Bw�i[ɍG&�-���>A��KH~��u���?P�����^�|��ս����u���}9.ˁ��S�߮,Y���b��W������z�!�oII�FE��_��I?-��lBX�]l/6����*-,%k�gg�%!�c���du}�*-BX��\�����{�~��N�x����'�����qI�:���U�[(�%�������$��
ܙ���?\��2�.(#U�6:�n�Cu�BN��6P��p���^�#h8�H?>#�{g�n�T+*(P�:׃��J�q�ã?�ǚ=�zV��$+���$P�ږכ�77��`����� ��x���v��X��F��M>]�T-���0}$O�8?R�"2�V1�]8��X=K핪w#���_q��+��V����Y����
���u����"��O�{��J8��5�X} ����n��S�,���O�{�J�8A����VJ5�س�1�%,�BKT�
�?�`�?���߿9���9獌��wMj��םʍ�J�U��DV��?��*�ƈf��O�� � /� ��@�ӭS����7*Dp�tG+Nc�0p���R�嫑�[��=l���2I�X u���D��Ш;�ٯ�	jș�q��fi_pz�/�����Ж ·d��N��{@_W�d����q@lddt\V~����I�UAc�߲��K�Ǭ�s%bL^�h{�2��E�gZ�2������L�pC�أVz���F�P/�7Z�����߃��;j�az�P��UH���2|�}V�^���W��F�Ǘӡ�z����j�0�-�y|�\.�V�:�X�����?�[A���8��C�s�JA������8 Iq[���=	���B�9럗w�O��F��w*H�	8�"�<KGW�u8	 �<��%�-
��*�OJgٽ��^�Q�:�K��*����2Na��k� �����g�0/�{#�B�
��XW���!;J���&�FՇ�D?p ]씳/|����qp��1�Bzpf����AB�Imֿ�s�0�u��A�L�<&�X4	� 
I�[����e��f�t�åtF?�f�"c�б��㽛;&�X���	E�
J֔��kz�/Z�py���`�%w�Ե���H���s0�H��BA$��NS�H�6�?�8U������|\-#�M��FwkC���SCϺ6%͒g���}�8��`A�����v�q�!�o(��J�F��%�h4z:.J�-D�-d
��j4�R��R$�S��0��l�	W��_>/��:⸑��]h�;��c�꽕d��]�,��E���5p�E�D�R��{٩�~:yH��6］��$��b̬��أ��jYbr\W�����|�|�i������9����[�˥L=qP��ʹ����Zά����B�U&܄�够��Á�JcW),JԳ��zY�n�
�E�8���q�*<OR5 �U���������o^��#g&��'�s�}����x䕊�ꤼ��hd"9)G7gl���"��v���1�%�����ug6o6))2cD��͵>�.�����\��A��%�_ߞjj�f���-/l���%��Q�a����~˃/c��!v�q� 0��7��u��O�|] u�՚�l%�TPh�� ,�o��Lr�~����܈]���8����"�a� [US�GE�s�B�-��� µà��������t�/�W�t��g��#��Z���rZ!�m_�TbFp�O�����R7���ԇ�D������ned�d9��ܳ��eqQ��9����ד67�����yh-O!��CG��@���j���x]ٔ��'��!�A�y�)��/�#��_�����~Y ���G
��aM�8Rܺ"߭�.ksm��2�y�� �e'9�q���^n�g�g�K6=Y�v���!�5Ү�f��(��'�.�_Cs+�������#���d�p�$?�B�<}1�?�>�壯`:}��?z��f[�&�+,Ȩ�Cc*��ۻ�J���?��"�G7���a�ÿ:Uɴ'U���U��\�M�뺍�Q�z����l�:|_yO����B�Ngy��iR��|�Zwlʍ�k�z�����~�e�N����f����2�=OZ(�b>c�cjԍW��"��l
��k;��!��d��s�b5��[�Z3�W��N�7�p����^�Y�`�a�g��SO#atͱh�5��R�Xm���9q;D�� ���ۓ�e\2��^H�KSPZ���3wER�/�/��h��w�������Y���"�_S�e������㩝+�OEzs��a�y18������J��Z[l�g��	�m�8��΍�54���ѵU�4�ӠD����^53�e�ړ�S^�kk޻1H��*��B��yO�X�c8�E�E��&5���l�T5�E���ei�Q�5CT��4,�k�kr���1�'1�Z�q�t�}k���\t2�1L�%��� ܨ8�粗Zr����wj���V�0��h0wr[b��u�b��i2�����.�6]#�[���}n��>y_�|B~Y������/�{;���3�c�O&Y6@�Tu?���Z)Ӓ�*1�]������8@#=cY$eߛp��;����m@U�\���O�
�c��e��$0�Y�0��;v�\T��j��<@dp:���\�&.+�[�A����x4�'�nz_%θ�q'��Ɉv"fN�ťIM�h<
r~H�ޒ�]�"�A�0�����J�f-{����6{:�,�nԶ������/�h�`�Q�Ch�%G��Z����-�(��B2e
v>-���M��j`D����SRd�#vS��`�{I�g�@[�i�&�K��^Ȫ���˹�=��d�B��͹A9��`s>���;���^E���Ik���AG�B�1�X�����ؠ������e����e�3��	��l�6�ߍ�̎N�hh���8+W�����;��ζ�f}G��I���c'����\���|�'���-�����B��ӝ�tʈ��	��L��"��gભ\��i�S}l�Tǖ�H�y�x���Q�3���'�%�e�?E�A¹8̌��PSZ啄�C�r�bK�G� ���_���ɂ�|��h�e��`c�%��Ꮨ45n �޽g�>cdSM���E��g��$a�S�K�}�3Ce)M�b�\8c��5v7d52 =v��JceU�)�����:c`�|�9�vy�/�|	j���!V;H�ek� �A���z8l�8;):�9zrT���5��Xd���DM{������A���#/{��2̫��"
��aq{�V�z�.[P� ���6Z�M:�~�O0" oIR�wFS�e?�Krz5��K�.�8É���*���A�ւR�3�#�$�,$���&���
�'U�H�f�_ae��D�W.���|��n�����tz�X�PYr:9_��r��-)ԭ���Yw��w��nS3��81%��R'6�~�)fG�$Tu�@�n���SY��_��HH���%����BIX[P^�g�i�n�E>}����F^�3���I��5k~Q�c	F)�xF||�aCH����k􁶱huS<&�~�d�H~���z`g	������z)�bV��Ɩ�ܴ��/��)�q��e��¹jS�F�I.W_�f��|�Րs��$��z��f���f�AÂ�̤�P��/*�;�BÙ�Q�������^(��f0�F�#9:����\��o�.<S��>����B��@G���C���%~�Z)D���Z�mE�ԩ,����Y�]����"��aĲIK$����y����֋����E�i�^�H��F����O&�?L��=Ѯ.Kr	-{���2>�.���:������.�?`I�5}�^$�����:�B`H��o ���e`?a~���CQM�@r����V6$i��^����젘zEq�M��H�
ۨ=G�YB����}hv�&�~t�9�Q���mx����O���}�>�i��"�7@o�ź%��3D���q PDOk#�A5�)f]�c�R+���TKn�-���|��vl> j%7pj��4
`L)t�y�
,� tU��	-3��G���X�n��\��{K��Ѽ"�J���٦J7��^W,$�-�L@˚] �H��t-=L@:�K�����,JJ�
��۞u�8�%��-^g�{͟2g�����h�d�~����ځrlm��G�^䅵�Z:[$��͢�@GlC�)2���4���A�߈�"��K2:��
c�.J���kD��YF���{�'��[��&�U��'��$�/�%k�?Ѫ���ܨ�=˻��{��yY��I����;�W��v�o�%�~$������P���
}���>[����:U�SH��0�	CL��Gv�� +�Q�z�_����տ��@�I�d�2�M>�h`��m����j3l5��E�~�q�x�����:���ܳ��s&��Z\����s������(gW�2������ey��s�^HM����aL��L�0�p�d�e3�`'n(IW�:=�����uJ����=�]�-O$KBvґ&떜aߴ�E�R.�����aH=X�V7���Z���Ӣ'�
=�7�#��H��UT�fnj7wK�;��'�ܠ�DEE�$}7�X(���s��u�W+�J�P�F�6$�Pj	QZ#由D���a�[�(�:|�?	P!4��T�w��mXa�#p;�A����v�e���RYN~\'��EL3v�ǉ*_4���0ꖡ��!���O
MjUGu�y{���?�Ә3+p�Z�S/<,c�%���艹�0�qQ�����'2���ʸ����#n�%u�Y���h��8�J�.�[Z��	n߾� >���ʠT�c �ܮ>M,���l�G�.�Y���OrK�:+'o�J,��uŦb�}XYj��-rx����}b�趟��Ż4�?��Z��\U�2��)n`r�����;,��Q�{�`;͡Y��i���/����G�N"?��"��1�Gt�O^;}w����F�����^E�.N�����xŊ*����¸��[hT~Dm;�$6HD��S�F0yۍ 3f�8ʙ#�J��D��%"Px퍹-�	�Kc��A� �Sa5埬�w|R���}��I��D��n�K�^�j���oM�:p��츍�]�~�N'���5���-�����܉����S8#��0g�7���׶;`��5���+y���ѨYT��X��z_�$�%C|`.9�ޮ���avͺG�m��
�i����:i�m��`jq�h�h~��#�0L5��2�Q�no�� ٮy/
l\\���W)�����B.��Bխ]���հ�%Oy�й|�F�
Gz�-
���t^
�j;-�*�@��e�f*���";xh( �f�q֪*P����w���;d�Y�xC����֥��/��a��gper烧gW��AJ���P\�+�Ȇ�Tނg�J�O�[�;`���c��~m{���+�/%����#��P�s�i3y{pĴT��FR a�<Φ��R"VI/�$���(��K,�J��Zyt�+�n�X��ɪɢ{������Y#�Ll��{؅Bf��[Á�!�.\����.q*m"[Ջ,�)__?���.���Ĝaj����nvM�^�+�'����T�5~���[�Q�_y�h�;c��<��
 zz�"L.���Ƞ�+�h�Ub�4��n�)��}8�xĄ��T��Gj���MQ	J·S��ҳ�H����?y��T�fr�"9�X�=��Zq���U/~��iP�[�j�Z^Й[bŌ���+A9���9�#Hv<9��k�{��!����1�h����ּ��?\h~�����x��'P�b��k9�|�V{@��:e[���b�P^�"E��x�]ͻ��X����V=>�4�hs�.J�w��j	�y�K[X�$L�b�o���/�+_)�
(���:#��XZ�aѸ�d'���U`���YZN�Q�Z��OY�N��o�ݰ#L��~�p/���������L�&M|4n;"�l�'v�/�\��dT Q@��>asw�o���}��f�Sĥl>��^������2:�v���S�u�����r��I����@�r�M��R���*����F����_��|�¬"����%'��~F0�)�@�+{�#}��,f�@t���d4�LI[Ot����$����9����b�x_�G��Y��P�FKZ�17�e���^Њ/�����-k���gN������n�9n�#���ݣݱ-JT$����6���d(��
�u�Jݙ�kև^����NT�u�Nr,����uN���zՇ�L<��/�t�{�������A�:_�t9�Cq�j~�S�,��u.���f�RJ�������{q��f!��^5� �)�$4
B9*�́��N��:�RV$�9��s ��M1u�1����ˁ�S36A��u����[���KWp7���9����>?�!ͭ
;[`�� v���@���|��GE}��I��˨�Q���L������Z�q�F%�tc�۪E�ᅗV�EOI���X��g�'�I�6�����=4=�D��3��ԊY��K'��[x���=ıQz�����TQi,�yF�'�$E�:�@�`��OǖrE_=�_3�Ud��i�`C�鉪OK�Q�x�t�~�x��KLL�ۏ�4��� ��Tpr������՞����{�ؑ,/y���_˘�b�$2sA"ڿ2���3O�(�F��	J0�	��)����4b�7&�Ѕ6��$�h���XP_�,�w��:~q�X��P)����"����X��I�W���yn�H���`񹹌:�������c������e�����*���.bG�0�vjkȪJ�6�R�'�N�Ǖ8|Cmc|�)֓B���;�"��Wׂ;�T$n��N�Ł#�f����žQC�tn��	dbX(�XJ'>mV�}�Cz��n�2 Z�ґ�
�e�vI�҂��/�I�䮥�Ha���u�,�'����3�B�W��ՐSY�sH���+���$��(����cc�>�o����f�P)�s�v�u!�a��>�[���H*���@A)X{�d�Bjʐ�Ǎ�.�BN�Cv�Ӿ�%C��`Q���@Q��Vk��3j5m�V�p����""(�b�c+���3֓���JDat�a���6�L��衩4���T�L�O2#ّ�y�ݯoC֕)���#�� �6k��(��f}�7��	��F�x�j�:�L��.
�ַR����$�0K@��n�9.�	$��H�B����QX*�TCӕ���a�?ل\���ѻr҇8f�1����u�(�]�����^�&d�H�ܪ�{��y���Vo�T�<��8t�JP�SV�&�D�_������c߉> "�14��Y�70
1��y=Y��m��z���%�^�dz km,ibt�W�lG�v��tbZ�ۑ���3��{-;Gw������X/�uR9��<�4%�UE����n��NrI���ǃetn#b:�[`�<�b$��ݗ�$�xV���@�댨8}７���|�z���|�����d�s,���''4��>�@�}�� ()����
�@p������%z��Rl`Q�]8����@����r���ր5����6�b������R�L��KoW�}k��-�.fy⇥�[@�(�g�VX�>x�ꓼ7��i��d�d׌���Xlʒ�і��L�Ҝ��}�z�3DJ��Ύ�`��P�9-	-v��4�Jg@Y��t��9���C����m��/�X�AY>�f�O>e�_D!�c I: ��/�wqn�q_O�=��M�62;���Y' /��h�;��% �C��]ס�|�Ct@���E<_Y8�Hg���=�C�	��歛(3�5&��L����L��&+��@����*��P	�]�ݍc��0(|&;{Xc�rt�e�2�?OZ[`ȫ`و� "ƚ^�P�}9t�s�ˋ"���c�ʂ�㸦�@�T�;�g-���jN˒UzsGG9[-�E�Qe��_FPӗ�#��R�T���4AĨ�Lt4�r8$K� ���JىB�ͳa����2�E���&���J�����⢏!��M�>$���$����U��i�DɊc���W�N�Hy��WG(�8TK%>v���;�Ͽ,���;
39z�^�a��͝�IO���Z��?&˅K	V�9��9.���Sp��zS�X��������c�����C�IK��`�c�tr8A`M��>"k����n�˂�~�eX�U��&�`�9�r�A�
(	I,Y�ɿ�Q�d�;�E���|�6��e�SN)]�� K�����)�iv�:{�������6n��-/��X�;Q2�ދt�T���o�u����S)u�i+($URs�(mɤ^��_6pg�X}����F�"�H�W�a,����o0�BA,���T$�b}	��+6V���۪4l U�-�u��^��ȬW|M�z8-?)P�f�`����S;�l�l��,�C�auN��pc��k�ͺ,�)�P������P�Mx݆4Ԭ�h!7��oEI�]X��"�O���^����b-[s��i:��+7i>8�P)#�3�����3H��4gȣ�oO��Px����l�S2�s�����nIj�mȷ`8K@��Z����E�[��gC�V�Yf.;�����B���T]W(��Ce���[>��Q>\��,	�ZJ���aʤ�h"�v��"�.5��}c�"C���3C˅.u0/#�y\9䞈��M1\������m�Cv��Rp�=tȏ�ѷ�����9I��Y�:�"h��Jx��$�O���?�ZD[���qf���}��>�WsQ*��/�c&���T�a\jD���\:hC�rcpn�f�do4�'�Sb�)N�/��	(�����?�\���ѽ��6���0��>�`��Lp p��3�<����!7������L�k#Fe�,Q��-<����HɩH�k4W"h�f,�����/�b+>�.�<#�P��Q�V���gaO���9v"4����B�˰�0j�.��m]�sccK�FV-����jSբXۏ�u��8�gV��E�.�E����.Pn.�*�*�NaRt�ryT/-FPqk���JDD4�ls(�*D���+�X�F ���M�ʰ���Q$ɸ�$O����Bb������ͱ�+�=^��?$t�l�Ͱw��M B�-�,�m�W�5�4@"����|�N��������
��>36�2��6�-�w���p�? "�Mz*"�  �q�+�1��I�A/|1_���v=M:z��ړ�D�c�ҶsjC9%���B:C�J�3����X�k�-: �5�q�P�c�QXT��NP.)㩝�̱3��F�h/��t��ip��|�Mbu���ډ�0������MVl�N���UK��K��ǅ�],���]����q	�6Oz��J�"p�(�mv7M�Wu [|�-4��Z�Yr.�	!<�\��ceT���]�Wq@�d 0j'���#���=M�_����*V-8��&X0�²�Sc�ї�,B�����$��%B����E4	g��Z�Q+�JV�!!�H!tY����/��� -��&�d�Z�>�"Z�&�s�F��ߨk��$^����p��R�Z�*��ӛH���W��%�v�_��Yڥ�)���WN_v�!K�$��Ij��C8Ml0:�W�)���>%���j|b�0�e�z/DyT񴐏��N0����q�+%�cS�'�����cA#!龈!��5���}5rך���.�~Amwc�y��IC�ڞxw���p$���S��� Vfgz��
xaj���Ż��v�8������0��E�ΥfWz��T:b�^�
&���jo��a��apE���͝ ��?���T&Yq�U����T�p��51HC͝��c������6�/��1:)EV(����8n8�q5�l*��>���ܩ�Mحn�;ˇ�C8�M��"�}-/RW'�x,hK��;ac�k����D�q���z�g�7\ͅvm{W�I��~K��b��+�R��m�7�dP>W>�Q�~_�;�Ou2EuAY���v���	3�	q�����3o��SO=�����N�&���a�C�K�2��爽�%�o <����I�$��@�&�貶���Ɩ^�f�C����1Q^ݓ�ʝ�����!�(�\W)���W�xmI��Ȫ�O��i�5��u���3�n�v�ف�}H�=��#���������a�������c��c�_E�-���m��T��p��������T�]uC��,�]Aԯ�/�!#����&�2R~���7.0⶟��[kr��D��<c�|b�fF��;SW��V^��"�M־t���x!p4�o�:dq��V�,�[��Z��=�H��f$i[��&<r�Ym^_��XR\���2�=�*�>A�T�x��a�u]YQ�'}�)3��ē�u�C;�a.;�
��T��_���le���NDL�5�[Hq HR.�AO9����)��]�6�n� ����I�Ͱ�>GK���E�=�>`�������(�d߯��ꓰEsta�֖�g7�RVd���kB�f�:��^��6���^{�Ĵ��nym��N8vz�F��fD��̠�&�L����F?�&�lk���2���9�P:A}�����jd�8��F����H�l�f�BQ�P��������({���Bc�:��G*�w�T���>�}��ˉ7�/��y�lm7�n�]Ƞ���IY��P��d��y+�W/n](���z@6�X�K_v��,��*V�t�%�E�e�	:�tp�|"�Q-a;�9���֞�x�])��C�A�v����A�aB�4RZwG�~r ��r+Hxkd��,ޱ�Z��/���!yuz��֚:L<6P�q����fP�߹�d���0
C�8�������l�ݸ���ZҸ���Z* ɵu����&bl�=NJw��4'��-^� �I�7��Y_��G��N�.K|4\�u]:�jo�Z�C�9�.*ҳ�dE�^l	��k��lF?^J번Q�@!wfD�W	�/=i
?D�MQb�zɊ�vt��|��4����1�n��l���o�,\�j��� ��сϯ��q"0�f9#���.�p��i�B���τ���� 5�.�ݲ���������V92]�æR-�ʷ,���A��N�8;)qS�~��+��2|��9״Q��kq� ��4)�,#>g�:��a�%����{�UY�<o����M{U�n�Z���{�X-!�f�j8_2���[��b�l�,����d�_��S�F��$�l�_�e_�/+}Xdp����mq�7,=|l4M;�Wh�';B��s��Q��R�����ȲM�c`@�t�ߊ&;��뫀m��1!|��S��e������@Ս��Q$�䋔��⦈M�]�UkLoC���c�������m?$�������)���Q�H+�sMlf���:��p(v�M�g��,�Gdg"��t&�,\/o�2h|+s��S����门��ƭQ;7 �O�eao5���9�`Ĺ��4�Y�
Fd{~��1�IC�5���@D^<�ʜu�ǡ'�&J
_�BЊC���җԫ�<�L��o�_Y�pbT�=��H6���fA�������#�?ljf�Mm�wdm�@��:�[��<H��=�?�gצ�Zۄp3��/~��f��+�+��A�CI-�0���I#Y��'|W����#;^Q�@6.W���_'�r/%L�Ēv�!�* �޹��L�f�j��1�	�_�f�I���t�v\�w-VF���E����+�H�ʚڟ<�T�$օ��x�!S��O�6��*��P�\���&E�K�u�$ jU]���ÐI�򮠲��_�1V��|�*�Q�7��g�(��l�-���}�UB��=)���A��B��8?O�a�z_t�ʏO�c��� Pi�x��
�]�ޘ�-�M�bl��Y�ث'{�Ȁ"��E�[՟��?�K��O������M���/�j䇼^
3��K�c�=���T�
6c/Ch#F_�ˍ�1�Qi��G( ��w�ܘ��B>I.R2-3��m|Vs1ee��K�df)��Z#��P@9���Zl���}�+R��4��?�S��ҳA>鸄7�k��E��A-9���>t��p��u����Cp��#ܒ�K��\4# ������}��(@Z�:���EB�Ϲ/	Q�t1�خ\�^<�#�1$Nuj�B,��K�B�5�G�b�_���kj���t[��RĐCD/���ʵIx\��ʓ�ʗ��i`3e[��c���h��K�ȣ?`,#��
3Z��R�VIQ��`&�3Z��G���=����K��yjůd�-�٤���xq_��ECѦ^G:�3(Rݻ$��ۓM��}G��s�׮z� �+p���t�t�|�qUȣD!x�"�6J�)Y6C0�cex�pH�T6��L���!Շ��=���}��&k�}���q��౸qTr��9.@香&�ǶJ�}��JN72tP��o�Ɔ{�jIs��qQ1W ��q�^P�Rj+�x`�brUs�MiƟ�zN�#�@�6+�i�Q�B�d�NO��A�a�٣�u�r���E�o6
{��1Nר�x�fZվ2��U��2D�"(��]26{u����J�j�{dr��<"��8ԮH�L� \wS���`�	��M��8��C�d�sKfJZ`��9��$��1�ֽ�?���q5o��K�7{����D� �#�ݪ(�o0����#Fb�2 �H�T�[��r�]XUqCo9Z�S	�y�R���D!ގ�>���?�
���*�/�_����6�ص�����-�O�ٽ��oE�sW����B�5l�j��'JGj�b�� p�=W�y�8z��Ii�a6V��9�R�y8M�� �$Mc4���ڸ���� P5��/���C�N�B�7D՞�(�L�2~��������;|�����o܇j�I�-��%9B�JE��]ܩ{�zk,��}gX��=kl�����U����򀹥n��?ר��#�o%M�D��TΣ��'g��A�Zp�(?�7b�)i�������>�j~3�8�r�g%<;͈\���V��m^�|4�]�g�&�
I�6��A9.���� ��L4js��e��PYAu ��l��ª�(7��>,�Z�?���Fq׃
O�Du� �B%�cم��ff������b#��d�S�Qm���T��Ǎ�SG_t��-<��pK�Z"���jR��H�?3����]Y�v!�m ���H~4hOg婚 ��k0"_Ϩ���&Rw�F���Y�aA��r�
N2e�d��%�.������o�R� �,�a�U[��<,ta�qC�l7�.z��z��A�0��*ӟM�K`�,iӗ\�<�N����-�F}�z$}V:�yh?�5��T )�g�5�U�v��f��{ a_o�v�+��;ף�D���/l@X����kA��D]�͹�J�O�K!א�j�&���6�Y2��m���6�A�{��;aalǅڑ���ѥ(�Ė.��~D
Y�,;וRU�-��R���r�"��~�<�=F8۟�WK�����Bi�����>��w�?,}0��~��k��F�m"��E�;��a�䏌�-m~��b�����4�4>#��S�q��M����b�`���dQ+f�j�d����^�7���;�w���&�,<��+)&;ʊ	Z�|�J<4�Z�!�mK�u���G	݌z���6:���[����o>��{L�#,Xh`���6������=�y�&����V�q.�Bl�l��b��ׄ�[s����,�0�O��h>ڋF�O_�%T�9��ײ-YfH(c�C���A�w����Ao�o5�����?�D���� �	�Ҧ[��a ����ӥ�^�ch��M�fz%�
t���p$T��	��V�p!��쵿@�R���Z�x�301�5�l��D�Lxfwjx��:{�g��ݲ���s� ���Ye~�zJ��w�k�֗sPa
>�*��$��b'e��
�6��2�������G��7�T�� �Ań�D��LD��Q���!�7�M'k𥼩�b1�P*��9��c�b:�>�(�3���nEy�����4Y�*X�Ij��w1[q+>���\���%4��W'�� )��~&�.v�}�#0jHeS���wd풷@�Ip�F���K�S���C������E��F�
:t�X����+	�ً4N��w]��6��p��+z���[M/D�Jb^)9�7��|���@B�:�#7���c���k�
�\�{vNb$.�$l%i�G8o6���^��OPXj��f)�Rd��g�0JP�h!J��rr�P�$0�+����N8bU�D�����,4/Y^<���~�59���n����E��)�`�a?��{�g��&Q?���f�Y_w7�"�,�������C�3�-m���f�naU���Ml7�c�!�yV�=�m�ĺm��y�/���Ҏ�S����~���N#�,(d�Q��pi�W^l�w	ȏ�3g ����J�C /�Y���4��L���^)��#䵱��􌰵O��)'q�8�k�|��$���C���ZT�և�1��	F��	q\�:�_�NUe�BL�}��]�5�2;�Ҝ�J(rL��������<7�Q�u��'��SH����VӃԞ�yƸm��G:������;K�!5�<K�E�:��Uײ�C���-�Q��k���_	v�tu��E�V��D���O?���D��I����T���ϖ��W� �E{h&�@�/�.��w�������ꔛL��i�4"ގ�R)�
$�\��r*T�jG&��-�������gD��	���-���3A������EQIk��&��Z���b��j�
����=��y�Y7�ZW_���u��i�A�j_���{��mf��'�l��n����1��6l�
��t@�O,ߎ(��="���<� e�C�����Y}�+m�j?B�,�7��웹�@��[������F�7�iE|����|޴0]-�TY���;� �)����gUoW��2�;J2ko �OP�I��ns��C[�}�٧7�U��_C�nUZG��AM���9�Y�I�A��\�U�,�I�3roTЌ>g��3኶��QwLqp14���&G����C2�	� �<T&�}���S'd���d������Q'��)���y�}��j�h�6�Ѧ��U�Jt�u��Έz8l� %\��F�J,�Ʒ����::���˺M�7�"��sG5b��8}iM�]}�ꧩ>+��.����+����/,���@��dZ̳�{mUN�k��o���{���$9-{�;��oM�I�u��Q/�0���NT؅�!wZ����q��+RWJgq�Gk^!s� w�R�X��NDxg����p?>��mG��4��s�����̄|
J������/�Y�QS�Y��ҹ�0�ߐ�����N,R���\��?*f�Qb�7��c�f����N�b�A���N��cc����o�o'Jf�&�@��8�9 ��% �y�Y|h;�UPs�fQ��N�HW�c?-#<�4�sf�Mt�x0ֳP@���~~��%֏�J�mΆU���1�ܴ@u�N���>�!�a�n���z�;d��Ȕ)�l&R��]��l03-~,�N�n3�lS`C����g8�y��V�i�{��
�+����]s6�t��d�g����<a�m���޶��n�
��"
��M����-NL.� ��� �ҔMp�j3qP@:`��D7�c?��(�����Zyxqt�=���.8����+ܖ�
g���%v��������BH[��XϹ�ER{��U�A�#�ՠ&:ںk��Ò� ���ߓ&��]�C���=�t�:�����b㔞�>����*s������yXe����@�y-�+$YT���)̕��X�/t���c ��M"���]|5��sD�:6����»m��Z�I�0���A�l]Rݿ¡R�<�}�XL���EO�d��c�ǚ�:oٖ����\
�xC�1��T�qpe��4�W70��1�
�#�� Z,�����X�w�S�ZO��U0��#�-q�K��0��	�� ���9��_��U��6������V�5����!�0a�]t!��B�j�ƱI��lj0�'
��c�,��!�@c(��X'a�_6:w$
�ۻ���v��~�H`�%&���y����OS�7]&�[�c͘q��m96�h�6ĸ�[2)߁:�����u�
����k�Lpc�%�+w<��PH�^��9̏�G���@`�N��@��d�3�x�T݇�"��,��l���n):���UX�s������-�s9y�/v�)�u��?������-������T���ST/�M=�	�$`7o�Ͷy=+GmGK������ъHQ����<�"��m{4�%��F����:��1+�_�\�s����%���l.��zY����\��qt�<A���%�ܛ���#����q���)�ut���ͤ:]Bƹ�zw��F���60�������?�޽o_CB��Ӌj6f�K��		�U����%�ʨ��<���3ZZ��H��`ZsaL��4IJJ!p섬�a4�s�~n�%r�D��w?����IÄ������C%�B��!��ɗ<5@�ȕ4��֟�����ݙ�����'�N��*�X��F���|*.�H�}B#m*ѩD�S�%,�1x��ܸ�G.K��8�Ϳ�tl��rTG���(/D\߬��u�옊%y��v�� �'�z?s2������;�+W���k�����.�������p�������W�qH 
��,}�!I$ �-Yn��ۮr��s��N��~m\��$S�Rh9�e��O��v"�`���T0�
3c��wXqjOt�а�!��:��X��j��n�s���Ϛ�����^����9�|_���L6�f=��4�[����e�@����uU+���,��ޒ���TF4���lFg�� ���_�֨���Kv�6��p�N\���xlc��nb�	RCu�e-ޚ<��[eP7{��z���_B�";v��Ӏ��D���8���0�O^ʶڐ;�^�B��eU.�Em��j�i�JU*���IZ<눻ݥ�[^�B��!v?��YeT��-SY�CP�M\�������X1S�K��EF	��z8w4&ngDI�R���A���<l��
;�=�@���-�<�[/u���
�d�N]�h��z,���GG3���@�}�zD��y�� ��Z�����G�G�gh�IMy��u�
��i �.�1�J��zi��:g��ˢJM���6���yc��%��õ@o� �ֱ��R�*�<�3��w(�`	h�SH+8���5��f��j����L.~���v >Ũ%�h^˷&;�yFY�І41��Ou�v�܁��Ik{(���Ƈr�>@'�a��#%@p���%g�wU�3�%���4O'�t��w�/$�����>�$��j�/��e��������РrE|��� �VN����v�h�0��~���J��`2�s͋i�B�p�Ԙ�4��i��U%$uU���-"蟼1d��y��#[�P.^��if��<�JM��Q����'��2y�;@`a0^���y��{��"
Ķ��^#nDO�T=�������;�'��X�4�N���%�& �!�DFJ�j�xdE?K�&�-�ۻ@��إ~9�k��C�4T��mP�N�׃�K@��5ǥX���cok��i��r_��l�nM�"�]�ה�%q3��@K��ϛeы��Ez�ꜥ�؞��]�y�@a���mˡ�5er��0u���Ս�)Zy�`��b�'�;�ۚ�t���n��	i�*�-������s!"�?�����u~m�k)Rv�V}^��}Zy��FW��cE0>--���BBV�[w�U��ָ��p��]	([�rgml���R���1욲u���t�H-�L�~�_�$w�t	C�=Y����6��ʶO'�MU�Kz_��E�yƋr�jKBsF�z� 'Oڍ�K��JH����a���8ov���1��-n�30��ǒP�n4I��f����a�� �zHv.�v3�e�Yao>%d�����B����j��;(�X�=i1��y[�y�ԧ�aen�7�X8�qo�K�+h�B>:�����.�I;��pl>l��M4J���#�cU�s�՘��\_�w�`�6�t����_�(4G�e& �4�7m,��!V��p�nt�W�܈� Dܪ�I�9PNգ�?�����ɨ5��U`a+��Njw�t�Q:<d�@�խ��u��6���8'f�Q�h� �Ĕ˓COi�D �ܑ��5∬9��7˿J\�>F��)]<�O]���W>��C6�ŭ>�����ݴ�Rh��!�D0���c|A�m�X������ @!Ξ̹�d�ǂm$���Upk�o�}F0��[P7>�� �J���a�or@�hu|SA"�<1�K;�zgx K0�0�?r
�>����NRM��:s����˿����y!�PPoGy�jx��pG�����"^x�o�41�j�����0a��.���;�+abT�i��o�7k�����f��A4Ui��C����R" �؎���o*�Rg̘�P��z�2Qu�Q�e�o���W�x@)����fKH�:��J_��?)�D�A�9O�+�B+�NE�����f"jL��EZ�4��Cp�nע����	��{�;�/�]M��U�E��a1����cwe�T1��/�9�d��@���@�jA^?	������UOp�m��{�%�ߧ���u���Y��R8r�Uy���D��i88�����W(����eQv�3p�8̮��c�	�?�x5���5a�̝z�<�	9敠������P�r"�S����D5%��-��.�}�X�q.��_��]���-y���ʘ�ۊ���5G�Q��W\PC?g�`b�n�Gqͫ�@)�\y�Io^.�$�Ex�{���~Ie����/�=^#]�N-?0��w"[�^��7t�����&D~�
��D�(]L����W�G��� �q��V!`�I�r�,��4˞�/�Ԃ���~�y�s�5ns�5E3��t�^�����zڨ�@���3Ur�"r�.�q�)@]�љ�<=�V��1봷/�/�$<W�����^_�ʗ���.N�z-ޡ���8G�p���O��$?��	��Cc�EG\��,�֚8�ko���5C⌼3�Lb���H@N�TGjZ�wQ��ٻ�
XS�?b�V!��
�n^L�%N���#��4!�;��0�o�>�orW�m�9'�2�>���aR�_[,;2Jhy9��s3��l���xï~̐A�H�U���l"�/{�����@�{�=F���ba�ٖ�ޗ�7�pD��=p0!������o�G���:iILO��ܛ�0���^v�滏1�8�V[d�7�xI��p�#%�[��/�l�=$���'Ϻ��B��O�
�đW���1�V��ځ��xƗ�%^� w����mM{�f�����]��aI�CǑ|�,;}֒�|M�1��cG�L�Y�hO����Zz3�	����}�e/xY��b�ܷ\*�^L�7cA�.3Nd���h�rH{�*�LR�����Jߙ�J�W��Q�K0�[9|�6J�IX4�0��2R-i�1 �4Q4����%$�m��xЄHl�z���]�ӂfk���a�7+������AX=t�5���)fHՓ���g�������Sy�;4��"&�����-w-����MF�Z�S;!+$r����|:�rm��|�O\�o?��j��̒���	�	#�S�M� ywB��(��/s$WL6���&-v9yZ`�D����G;�s����+cC6-�8j|�k]��I�g~<��D�3i�4��7��@>�:'처�����UrJ���U�m!)�܀��Gg��܏c����� T!�����>�g�����")�L�b6Cv���6V��������V�HU65h��C���}��@:ĠD1m`��\̼�1^#�j��K+RV��?6%���)`�E:1a0�1sAFb��?:_��4��0�<r�K(�r��"�Ew�*��%h	 ��3�jE-�0� +BΌ=Go�E�q�,W��G�k	�m�P2���*����a?��i�T�l	�u�A�7SϚ+Ô���_�E��uwáV��"���X|(l�gI��?T��}������2-�.�"Y�ϝu�a8�o������h��F���L��L���N��	'��j�շ��R]�8x���y��υ�5�����7B8��\h_����M&��i&��aπŤ����9��琥�ㄏ�xˢ��z��<z�DB��1�{�ZBʤ�09�5�R�� �𲁶=ےi�k�"ۜ�1���	j��� �u�a_m����mj��3�3fޣ�};C�#gx�aٜێ�"Z%d�m��~��@8?9�g�+�-�����x/���H�:�-�jƝ аČ���Ʀ}%.Yt"	��K|���O�x�=H��Ll���Bǽ��,�}��sՙ��V���98֊@�	��%�e��&7A�R��.<7�
x�~#�U���sG<���z`�����0^��̘�ܠ¡oE#��>�r�/�3��1����i��7Z@��������y@7��Z�U�^����+R�1�3'�]�ˠ��%_���K���}1�Oc�QekMB�:p^4����7�:U�ɚx���)�Y�/��居d=8���K�� �:�����_��
+F���H��}��O��Uϕ�� ����=����7Do?�(;��(�xO$a���U���!� ௙s���I��VD��:j/��%���n�d���N3[�!�W���/�GQȏ$%\�����b���V��|�T�Tri�de�}ɥ���ڷ���z]���0@\�����_�1�K�?������ʝ	�ܽh;R�iW#��A�تW��H����?� \��}R�8a�9�z��2̸JbW�mÀ�}���Q�pM�z���>P͢EDF�by��R�C(�>�r�(���,*���6h����B�F��>�X�-,a)gY�j-Gd�$�V� (�\���r��h#�����{�%�z^��W�wO��l�al�y��UZ�A�qc2��􊺕rn�!)^щP7��(���l6���Ii]AJ4n�)G�.[U��,���}����ڶ��q���X@��k�1��e*����g�ѫ���"�b�x,	6 UFM'c�D`溧��&p%�R�;���@� �s�
�٬c��v����톄ճ\��*�����t�_�;��d���xD�
n�\�z@]�K?��o��[�M�5���AGe�ѲR8�#��w�ۇ����ń�#�]Mbk��P�g��"�-��;�������q}#�MDڧ�k�G�M��0�!k�?�����f�`u� ��X�0@����¸=
�X�^���'�;/��=v��葷�T�2!{��-9�ta�.�S�_��������#j	����8L�Z�a�yq��0�(�jp���z�K����Q�E���GA#R'6��/��}3�U{�<��w�_�1�k��%p�`/���y����
~���T�?Q��;du�+td�|$V��Q��s���Z<y�9]ؽb���K���(kT�Gv�b�򙬐(Ow��Wm%�E�0O��
�21n�:Q���;����_�bQI��Q����U����{�R�5C��8�3���b��B"���cv�$+��&��ztʯ�//�������m�Ml��R$	�Iٲ�ɥ�G�QZ�x�|���7��="�Up� b9�+�#~�ങ�C���$%�q����
���
�hV�h��7���dpv��0��)��tB��a��_{����Z�@���M`V�:p��˼d�nʤ ��W$5�w�V�-�1���4 ���颊����9�Hӟ���L;��҉M��d��x��V��8WV K���Z�Ϛ[G��)\k��͏��iV������3�������B�!��~�ښ>�(��KP/OB��r�k�1얱> I*#��j��5��W�{����q���昮]�i��K�e{�S�C��BZ+���3ǚ�[�)n�Uqc��WӸ�$��oq��c�l�L�C�DVj�q&���+Vz(��[7OY����O2z;Qx5  	wD�iq��qyQ�Ý�v�ۯ�8�w^=ڳ����E��M(�ʉےԓ9ЩM���_�H�dX�|܃�Ӄ5Sb��8��% c��� ��*�D�L�b�He��F�-E��y����0{�N�,�|�u1�n~��~������	�承���*¶�*��  �9Ԣ���Cn�y`��[�Է[��)&�}+��;���������-�y����2\��EZIq�4�=��Y~�,Y��DgmQz����]�r?9pZ4#"|��#؛H��[ޠu�:G�uU6]s��c��Wկ��|HA-S:��uD)�`7��`��G�:�'.����"�`���K�י���:��w�����W�@���ɡ"�zh!����]�J��t��a�'�*B���dXpN~�>���*�>��M5 _F��F�m�M;����%��(�������|`r�j�:��2�/� ����ݚ-�Z'���M��ڟU��c�cB��z���?��>M)l���^ލp�*ij�څ��՚��#7b
�"6t k�֌)�Kn���k4�o���f`/ 2Z�n�Jz��Кsa�eAv�M��c����F�4)��Zhp�sA@o.��(�J���s���\��\�h0���`v�n��b�'�4n%�krC=��]�M����BOuF��\�F	��h��A�6�`�s��k 1�p�7;��ВW4��REh�BPⷔ��ޮ��i�_����vLK��L,��Vܪ�j��A�D�j/�Օ̺$�ݔ��z��O�J[e�D"���#��o߀8�7⏼O�.>,�~��������2	ƾ���!�F�\�Dk������	�dv~J�ͤ��ܺ2��5��g'g;x��
�<�L@�]9�[��gY!LsC��ʰ� W��;~`ה��(N�������Pv~�e���q�=Bu/�v��(&IwM{>ܽ���,'�8����	U8	ui ��_�-�|��TN,���$@W��@��=�{D|�QV�����ܐ�r��m�����h��������8G?*��N�7b'�����2.�ē���%��Gj}�e�79)f�Ϯӻ*31� ��j�~���qT'V�" ��݇�AG��˂�0伈~��g�/���O��Z$?���S�i�Z�'���s�4�9я������E�۬�tGS5�F���T����5.?��D�i���楄%�{�<��w��j,��~�a16G��z�1;w�܃k����_�&v�< �E��6Ԃ��D��pn�]*�Q��È�uؾ��k�!�4;NM ���5��ج�"�Mc��IӘ��ĺ:�P�%��>�D�0�cЏ��Q�L�Z4��bؖ1�����b!
\��ES�nz���8�{;��*��!��j��wy��)��d�8G�o�h�4��`�:��Wuq�9��,qCP��ܺ.t��&�~�*S�g��V[b럔���ԪAi��8dI��1���G�bH����2ӑY�!w�v��� ��_X��E�\=	Pځɍ͞0qDj^�Ĩ���Ua�{����{n&Zp�{9ud�J#�:}B{�� �ȅ�;NĜr&���b��	���*��!T&���[X��A�y&7Zk%�뺂���ja*ֹOX(��=����k�s�cs!�p1�QW��������*���
��b����ȇ2��Нy�+b𼌑�^�-v__�v˒"����60�c_�b�/_�)޸ ��E#m�Ds�%ioGQ|�6HL0�SA
���`�o���� �b�MG��`I����­p����=J��9N�w�K;j��BW;j��SDW�I�p
���g��x�ק�?oO������e(Y��m�e�<�PbV>�*�w�����u\\I]������~��`�E�%�ȯ[��C�#������`շ0<0�h/��������g�%]� Iۖv�r5��tx��9U�8n������#O��1ˁ?2�h���SLt���J}�u.��r�<��̩��z�l��T�<q��~N�/
P|PQ\�+(��>�|^z+����C=
c&4�(���@�36>n��8Ã�QZ�f��OO@���F�E��pr=0�<���잢V��"<2���I�~�D�����L�e8F}�Q&M/h:Qt�r?D�D��$�n�
E|'T�� �ݣC�L�*xؚ���rj��'el\j��;�b���m(�q�`��Y�? �tG��������‎��В�C¨��(u�Cg>&�{��#C�tE	R��y�*�ʬw=�_0��XKߺ7�7I��ꧠ���a����gfA�qlͤ���&O	�1��j���ذ>�XyIIp����G98��5�UU��I
,53h�8��=���)n��tj���j����R�~9���'2]��+�E@��U�	R".�����S*�&Q�'�#���"��ə�n�SU��4��6�N��U\Pѿ6�Z�A!��,^�������_%:����yS�i�zE��8�p�"2����̑N[ծ��{��j�D3w�^�8)^T��Tvt�I���R�8'1��~��l��@{����
���S�4g�c����$��"q8�^�I<%l�$d�+�W�]�[���KJ5\�p�>�6����	�^[�޻�m_����3vyו��Tf��_+���z���/�
�b��Vk�R�>��?��I)K�WZ71�����p��$��ZH�` �:t�+'��d��v<,�Nz$CX��D���;��Y�\�7eX�����$*j����3₈H>�Y"�&��n탸�q��)�j����άp�FL����$R�E���!�-Q/6���	L�B�y���L"9�?�_jE�Q��>YE�������T"��*��Qc��H	��_���LN%��:Lo^*��#�09C��q���i)�y��7��;�Y?g���ϻ���g�X��k��"Л�3ʢ��Ԁ�MJ^��Hگ�9�iP�*�g.�y�-�	km����.b�Hp$
�x~B��1�6� 5��
դ�oݨ�\�.�;0�,
���<����� �&U�����V�]׺#�����N�^��H��L��3��}���u�i$nI$z^�	f��v���ϙ�cbH:ת���k����Ξ) ����N�%�.Q he��p^pg`�����[�H0V��@KTD늂Z;��#�j[����ζ,6��X/-V�E���X�� �X���P��$�p��&ϡ�=t�Fg
f��x���=�C��H=�JWp����< #�C�A��������1�TO��(_���[a���l�S�nV���5Z1���π��iYO�3z*��nX�Ҿ��W6��vH9��|S2(Cj_��;M��:Y��6��ox�̠P���ph�ibw5�.?vh'2��&�r�S��{�\�I�/xyl,��W8B�c�V�̈́*ԼkS[ ^�C�������e���4a��g锛�6q�n�g؊4�wZY���~`~I����'�$�r�qØ�����f+"���#ڔ���w�b�����wdz�ܺ�w��>������U�z�"�k����I-����)����t�)�8���P�Y�.G�t3���v#����B��p(���%b�,m�����ڴȖ��'�Ʈb��H���~������\�,;�9}��Vbln�=i������C��:x�@��O}�6nzQR;Z������V�ޕ؉0U2T�&qJ���:�ȱ��/���	���vָJ�-%�Y*H�ɰ��/����g�yG�*U�E�nb��UeX�V�)	�R�O�� m�Ԝ��%.?�XdX$)������=:lg{v�_
"gH�A5��峔<>h1|�k�^������e��
��=�ȇ*�|In�?WVjH֐؈e\ZE˷��CY�B���Ss-?�P;*g��!UP'�����e�~eX�]�����|%���yL��ߪ�Ҙ�@��g���}G`&�b� �	����^nYm?�4�ǆ��`9w�4%oG���Y2$� !+V.�+����]7���I��G��o�Tw�!N����i�6�(�Tce\�ҍTC���1X�\�`�6>b�^�~�N�� ����иX�#I�q�}�ج�v�|�C�öF�J���oVE|�a��x:�c���;!{�c��,�ym��N4���^DzՐB����ee�-�J1�q�.�XD�s��+ �}�����F�K�spfv	[����5��c��]�,�����%C��Q����/����������u��,l�p��� Q)��ns�����b�sj *M�zz��IhGth�a�;t����C�<�]�Ɂ����u
@%�Wo�m;<��rڬSh0�H�k��?gD�J�[%��8�\	��s�&��zm<�v��s�V�������@��8���&��X�*�v���j]<�MI���I�+�4��e�g��e�/]0�,��tݤ�(º��n0���w��h�B�����I�(����/'�˘<��� ��cӰ���V���aъ���ȳ����jmyKM!S.IjW��Ti�<#���a���r\X�n~���_�b��iP����`(U�+��d��!�"@��N.�W7$�������;OŚ�
�Ck	{�"qpE��J��&��R�S��8�9����5P�W>"�(;j �e�s�����e�"�i~��%��NVǟ��0(�~JוPsl�6K����VzҾ�>
8���*��Na� w�?��{��d�(��v����Uɶ���*�Mq�h0��0�s�j�kszC�� �T�.���=�5�{�b"5w^��b�~�O��p�qb���gڒPg=�F䚦[�6~|P�p��J�v���E��jJ^Z��7F�F@;U�;�d6`T0OՁs��'IzjR�p	Z�c�&�g�cs~}��gi�vyh��Bb��d���$sqX��0
%����6�إ���3#�����ai?O�D�*�]����3������UqsF���?��"�s���r��A&��i̔��7x�Ҝ69k&#�v�F"@p���G`n�wؿT���ϖ�ۻ�	�M0�8%*�$�q�¹�Ӈ���ƿ9�Öѱ���aP!�ڤH�lh�z�;؍M0��Di�F��Tp��U����X��c�,-���8}n�1�HGKp!���7g�����i�X���r�W��V@k�`f�Q��_�ӊ���ؔJJz��+��c�f�����*�Z�!����ya���n�0���x��?��?�o}k���z��8�M�Y�!{X#f����Ç�� �j��:?#t���g��PM����p1�O��E�O�MzHO+=�쉥W��Ҵ`ni�o�a'ka@�>.��($U�S�fsa�Ϛ%N#Ԓ4.��W=�u�;?JB��./�� O�5��&P³F71�غ���N�T6��*=����/��:��2L��4A�=IШ�=�����ENs,Nc��n�\�^�D1��������'�pZ�)�+�:���O>�5�V��i%�r�L��6��X�W�XT/$�MK�@���Ԡ+(���@��_�v�BCF6��ؕ�)�zW#T���d+�yY�Fx�|B��U]��.A{C�*;T����JT�8�<BN!|�m�Y��}D�g�#V���Y!dFT���n��$��f������$�=i�ω�I�(�U��
���[����Yv�\$��[���;ߘ�N
�e I5�Y��H��đ�pL��l}�pG#��ܿPӖ�Z
$ȭ�,Q�zF�uI<��Af(g0b����f�5�gD�Z���i��!���ͪ'j�d�r�n.�}�:���af�h랬JS��g<ۏ�P�ȂTE|�1E�~�M��ew�z�22,1^3�a�Y��U���1�2���|��w8_h�j�R�#�Xخ� 5>z����������# $1��!2��3�	h\3����1!�v��F(��=+�[�X_�V.m��N�l�¬;h���~�E�����|A���{C��6�b[y:ۚ����3c��4~k���WH�^��������0g��d�6��7��j)��.pD�-�1�Y�-DLD�v� T�N��~��n�Ȏ�8�!�Ī��:�s��!Xj;�~2���X0��)d%DG�ֿu'`\x�zѓ]���w�Z��J���K0+�.,@O��yf�ȏŚ4Ǌ�P�� �c���j�٬N��R�׵@��jS����-�P�y��}�3-~���5�� �{zT~�y��s���P�P�V	b���o�qK�`3�C�m�&���׋e�y�x���S�`\17k�u�;��p��qע��)A&�I�|�<��E�~���]�ɼ����Uh]se��e,	V��{�p8z�<�_��*�B'L-��,75��PQ:��	WMW����Z^��8����Zk��cX�m���_-��"�r��>�sH�r1F�ȩ�����"�NL��L�C��H^��4!�>-عb.�C�V�Ď���,�	?V�w�n�O�\/]�3M(��W�~�w�M�t�h��z���.ϳ���aAwh\y�&��+ �,I]��L�VR�1R��[[Pɑ����,@a��FX&م�n�������G,n���W�2P��ց��|�-MI��|�;�ּ��Ug�imƋє
�柏�!S�\��H� �U����S��-����ߢmp<�oā��=Q�~���L�~�yۯtFw����Ҭirc�^j��{`�	pp,�c���Ql�Q��O�]���0�g�v	��.~xs��H�%i	F�܄O�B7X]�7-N�jŜ��?3p����F(@7r���b5�u�b���u�u��x����h����E�5Oq�J����x\ӄjӕԅ�6$Z"jVH��!���e�$��8����#'��������ua�	��*�$�o�9��MRX��x0�  ���CQL���ZeH�b��/?s�:h���:���Z}��A[G?�ͮ�(]��,��ђ�^���P��:���	N�w�"ރ��r��(˪���:�Z���'�5!3.̪�L��;�~C�Eڤ��F�Lշ��&�ن��ܲ4�Or��O&W�/l�4"&3؆�=�U���R�͋�P���+,ҳ��&��\=*K]@V�P�����+R~{}���l.�o0�Y{^z�������m�F�ϵ��Pp����~j'�u���%���������J��@�=��z,w,f�B@1�%�N�h�o��-|��ck (��r�6bW��[a��ƀ|6����JFΡ"S��6�oa~],����>dU�c��qΞtm���Х͓Z@�&r;aG�/d�-����+�p>��6h;���h���|���(��X�S0�KFX��/��}���=�pE�ʒ5D���ˍ@�tv�����>,VZX��V���åB�E���q��,�S��٘�=3*3��A��R_�47�������o���c.Ѝ`�;��mC���|������Õb��˭�2�%4�=Ue��ڸ�ǡ%fY